// Note: The purpose of this module is to convert the edge-sensitive 4 phase
// handshake input to a single-cycle pulse

module reader #(
    //parameters here
) (
    input logic clk,
    nrst,  //clock and negative-edge reset

    // Data inputs (received from chip pins)
    input logic [7:0] input_byte,
    input logic is_key,
    input logic reset_hash,

    // Handshake Management Inputs (received from chip pins)
    input logic input_request,
    input logic output_acknowledge,

    // FSM State (received from fsm state block)
    input logic [1:0] fsm_state,

    // Signals sent to the data router
    output logic [7:0] input_byte_pulsed,  // This is the input byte that *gets pulsed*
    output logic is_key_pulsed,
    output logic input_byte_pulse,  // This is the pulse used to communicate the 2 outputs above ^^^

    // Signal sent to the hash generator
    output logic reset_hash_pulse
);
  //module code here
  // assign a = clk && nrst; (example)

endmodule
