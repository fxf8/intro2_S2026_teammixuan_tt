VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO stoplight_example
  CLASS BLOCK ;
  FOREIGN stoplight_example ;
  ORIGIN 0.000 0.000 ;
  SIZE 160.000 BY 100.000 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 21.580 2.480 23.180 95.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 60.450 2.480 62.050 95.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 99.320 2.480 100.920 95.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 138.190 2.480 139.790 95.440 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 18.280 2.480 19.880 95.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 57.150 2.480 58.750 95.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 96.020 2.480 97.620 95.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 134.890 2.480 136.490 95.440 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 2.000 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 2.000 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 2.000 ;
    END
  END rst_n
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 70.930 98.000 71.210 100.000 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 0.000 10.030 2.000 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 0.000 6.810 2.000 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 2.000 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 2.000 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 2.000 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 2.000 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 2.000 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 2.000 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 2.000 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 2.000 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 2.000 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 2.000 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 2.000 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 0.000 3.590 2.000 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 2.000 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 2.000 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 0.000 93.750 2.000 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 2.000 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 98.000 61.550 100.000 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 98.000 67.990 100.000 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 2.000 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.840 2.000 92.440 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 2.000 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 2.000 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 0.000 100.190 2.000 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 98.000 51.890 100.000 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 2.000 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 158.000 71.440 160.000 72.040 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 2.000 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 2.000 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 98.000 84.090 100.000 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 80.590 98.000 80.870 100.000 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 87.030 98.000 87.310 100.000 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 74.150 98.000 74.430 100.000 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 98.000 113.070 100.000 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 98.000 64.770 100.000 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 0.000 90.530 2.000 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 2.000 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 2.000 ;
    END
  END uo_out[7]
  OBS
      LAYER nwell ;
        RECT 2.570 2.635 157.050 95.285 ;
      LAYER li1 ;
        RECT 2.760 2.635 156.860 95.285 ;
      LAYER met1 ;
        RECT 2.760 2.080 156.860 95.440 ;
      LAYER met2 ;
        RECT 4.230 97.720 51.330 98.330 ;
        RECT 52.170 97.720 60.990 98.330 ;
        RECT 61.830 97.720 64.210 98.330 ;
        RECT 65.050 97.720 67.430 98.330 ;
        RECT 68.270 97.720 70.650 98.330 ;
        RECT 71.490 97.720 73.870 98.330 ;
        RECT 74.710 97.720 80.310 98.330 ;
        RECT 81.150 97.720 83.530 98.330 ;
        RECT 84.370 97.720 86.750 98.330 ;
        RECT 87.590 97.720 112.510 98.330 ;
        RECT 113.350 97.720 155.390 98.330 ;
        RECT 4.230 2.280 155.390 97.720 ;
        RECT 4.230 2.000 6.250 2.280 ;
        RECT 7.090 2.000 9.470 2.280 ;
        RECT 10.310 2.000 12.690 2.280 ;
        RECT 13.530 2.000 15.910 2.280 ;
        RECT 16.750 2.000 19.130 2.280 ;
        RECT 19.970 2.000 22.350 2.280 ;
        RECT 23.190 2.000 25.570 2.280 ;
        RECT 26.410 2.000 28.790 2.280 ;
        RECT 29.630 2.000 32.010 2.280 ;
        RECT 32.850 2.000 35.230 2.280 ;
        RECT 36.070 2.000 38.450 2.280 ;
        RECT 39.290 2.000 41.670 2.280 ;
        RECT 42.510 2.000 44.890 2.280 ;
        RECT 45.730 2.000 48.110 2.280 ;
        RECT 48.950 2.000 51.330 2.280 ;
        RECT 52.170 2.000 54.550 2.280 ;
        RECT 55.390 2.000 57.770 2.280 ;
        RECT 58.610 2.000 60.990 2.280 ;
        RECT 61.830 2.000 64.210 2.280 ;
        RECT 65.050 2.000 67.430 2.280 ;
        RECT 68.270 2.000 70.650 2.280 ;
        RECT 71.490 2.000 73.870 2.280 ;
        RECT 74.710 2.000 77.090 2.280 ;
        RECT 77.930 2.000 80.310 2.280 ;
        RECT 81.150 2.000 83.530 2.280 ;
        RECT 84.370 2.000 86.750 2.280 ;
        RECT 87.590 2.000 89.970 2.280 ;
        RECT 90.810 2.000 93.190 2.280 ;
        RECT 94.030 2.000 99.630 2.280 ;
        RECT 100.470 2.000 155.390 2.280 ;
      LAYER met3 ;
        RECT 2.000 92.840 158.000 95.365 ;
        RECT 2.400 91.440 158.000 92.840 ;
        RECT 2.000 72.440 158.000 91.440 ;
        RECT 2.000 71.040 157.600 72.440 ;
        RECT 2.000 2.555 158.000 71.040 ;
  END
END stoplight_example
END LIBRARY

