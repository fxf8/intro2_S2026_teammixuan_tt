magic
tech sky130A
magscale 1 2
timestamp 1769113952
<< viali >>
rect 14749 18921 14783 18955
rect 17969 18921 18003 18955
rect 10425 18785 10459 18819
rect 12357 18785 12391 18819
rect 13001 18785 13035 18819
rect 13645 18785 13679 18819
rect 14289 18785 14323 18819
rect 14933 18785 14967 18819
rect 17141 18785 17175 18819
rect 17785 18785 17819 18819
rect 18153 18785 18187 18819
rect 22661 18785 22695 18819
rect 15853 18717 15887 18751
rect 16681 18717 16715 18751
rect 17693 18717 17727 18751
rect 18705 18649 18739 18683
rect 857 18581 891 18615
rect 14473 18581 14507 18615
rect 15209 18581 15243 18615
rect 16129 18581 16163 18615
rect 18245 18581 18279 18615
rect 15301 18377 15335 18411
rect 17279 18377 17313 18411
rect 17417 18377 17451 18411
rect 18061 18377 18095 18411
rect 13829 18241 13863 18275
rect 15485 18241 15519 18275
rect 17509 18241 17543 18275
rect 13553 18173 13587 18207
rect 15853 18173 15887 18207
rect 17417 18173 17451 18207
rect 17877 18173 17911 18207
rect 17785 18037 17819 18071
rect 16129 17833 16163 17867
rect 14105 17765 14139 17799
rect 14933 17765 14967 17799
rect 16589 17765 16623 17799
rect 14473 17697 14507 17731
rect 14657 17697 14691 17731
rect 14841 17697 14875 17731
rect 15025 17697 15059 17731
rect 16497 17697 16531 17731
rect 17233 17697 17267 17731
rect 19257 17697 19291 17731
rect 12265 17629 12299 17663
rect 12541 17629 12575 17663
rect 14289 17629 14323 17663
rect 14381 17629 14415 17663
rect 15301 17629 15335 17663
rect 15853 17629 15887 17663
rect 16681 17629 16715 17663
rect 16957 17629 16991 17663
rect 18981 17629 19015 17663
rect 15209 17561 15243 17595
rect 17509 17561 17543 17595
rect 14013 17493 14047 17527
rect 14289 17493 14323 17527
rect 17049 17493 17083 17527
rect 17417 17493 17451 17527
rect 16773 17289 16807 17323
rect 16865 17289 16899 17323
rect 17601 17289 17635 17323
rect 17785 17289 17819 17323
rect 15025 17153 15059 17187
rect 15301 17153 15335 17187
rect 17417 17153 17451 17187
rect 13737 17085 13771 17119
rect 14013 17085 14047 17119
rect 14933 17085 14967 17119
rect 18153 17085 18187 17119
rect 18521 17085 18555 17119
rect 12817 17017 12851 17051
rect 18337 17017 18371 17051
rect 13829 16949 13863 16983
rect 14197 16949 14231 16983
rect 14841 16949 14875 16983
rect 17785 16949 17819 16983
rect 15025 16745 15059 16779
rect 14473 16677 14507 16711
rect 16221 16677 16255 16711
rect 19257 16677 19291 16711
rect 14565 16609 14599 16643
rect 14841 16609 14875 16643
rect 14933 16609 14967 16643
rect 15301 16609 15335 16643
rect 15485 16609 15519 16643
rect 15577 16609 15611 16643
rect 16497 16609 16531 16643
rect 16865 16609 16899 16643
rect 17049 16609 17083 16643
rect 17233 16609 17267 16643
rect 19165 16609 19199 16643
rect 12725 16541 12759 16575
rect 17417 16541 17451 16575
rect 18889 16541 18923 16575
rect 16589 16473 16623 16507
rect 17141 16473 17175 16507
rect 20545 16473 20579 16507
rect 15209 16405 15243 16439
rect 16681 16405 16715 16439
rect 16773 16405 16807 16439
rect 12909 16201 12943 16235
rect 15485 16201 15519 16235
rect 18337 16201 18371 16235
rect 13921 16065 13955 16099
rect 13277 15997 13311 16031
rect 13737 15997 13771 16031
rect 13829 15997 13863 16031
rect 14013 15997 14047 16031
rect 16865 15997 16899 16031
rect 17141 15997 17175 16031
rect 17969 15997 18003 16031
rect 16773 15929 16807 15963
rect 16957 15929 16991 15963
rect 18321 15929 18355 15963
rect 18521 15929 18555 15963
rect 12725 15861 12759 15895
rect 12909 15861 12943 15895
rect 13553 15861 13587 15895
rect 17325 15861 17359 15895
rect 17417 15861 17451 15895
rect 18153 15861 18187 15895
rect 14013 15657 14047 15691
rect 14473 15657 14507 15691
rect 15209 15657 15243 15691
rect 19349 15657 19383 15691
rect 12541 15589 12575 15623
rect 14657 15589 14691 15623
rect 15853 15589 15887 15623
rect 16773 15589 16807 15623
rect 14289 15521 14323 15555
rect 14381 15521 14415 15555
rect 14749 15521 14783 15555
rect 14933 15521 14967 15555
rect 15025 15521 15059 15555
rect 15761 15521 15795 15555
rect 15945 15521 15979 15555
rect 16497 15521 16531 15555
rect 16589 15521 16623 15555
rect 16865 15521 16899 15555
rect 17049 15521 17083 15555
rect 17141 15521 17175 15555
rect 17233 15521 17267 15555
rect 12265 15453 12299 15487
rect 14105 15453 14139 15487
rect 17509 15453 17543 15487
rect 17601 15453 17635 15487
rect 17877 15453 17911 15487
rect 16313 15385 16347 15419
rect 14749 15317 14783 15351
rect 16773 15317 16807 15351
rect 15761 15113 15795 15147
rect 16405 15113 16439 15147
rect 16589 15113 16623 15147
rect 17509 15113 17543 15147
rect 17693 15113 17727 15147
rect 15577 15045 15611 15079
rect 17141 15045 17175 15079
rect 15117 14977 15151 15011
rect 15301 14977 15335 15011
rect 12357 14909 12391 14943
rect 12541 14909 12575 14943
rect 12633 14909 12667 14943
rect 12725 14909 12759 14943
rect 12909 14909 12943 14943
rect 13001 14909 13035 14943
rect 13093 14909 13127 14943
rect 13553 14909 13587 14943
rect 13645 14909 13679 14943
rect 13921 14909 13955 14943
rect 14749 14909 14783 14943
rect 15209 14909 15243 14943
rect 15393 14909 15427 14943
rect 16865 14909 16899 14943
rect 17049 14909 17083 14943
rect 14197 14841 14231 14875
rect 15729 14841 15763 14875
rect 15945 14841 15979 14875
rect 16773 14841 16807 14875
rect 17509 14841 17543 14875
rect 12633 14773 12667 14807
rect 13369 14773 13403 14807
rect 13737 14773 13771 14807
rect 13921 14773 13955 14807
rect 14933 14773 14967 14807
rect 16589 14773 16623 14807
rect 16957 14773 16991 14807
rect 14473 14569 14507 14603
rect 14775 14569 14809 14603
rect 18245 14569 18279 14603
rect 18521 14569 18555 14603
rect 13001 14501 13035 14535
rect 14565 14501 14599 14535
rect 12725 14433 12759 14467
rect 18429 14433 18463 14467
rect 16497 14365 16531 14399
rect 16773 14365 16807 14399
rect 31033 14297 31067 14331
rect 14749 14229 14783 14263
rect 14933 14229 14967 14263
rect 13553 14025 13587 14059
rect 16773 14025 16807 14059
rect 16957 14025 16991 14059
rect 15025 13889 15059 13923
rect 15301 13889 15335 13923
rect 17233 13821 17267 13855
rect 17417 13821 17451 13855
rect 17601 13821 17635 13855
rect 16941 13753 16975 13787
rect 17141 13753 17175 13787
rect 17049 969 17083 1003
rect 7205 765 7239 799
rect 9137 765 9171 799
rect 11713 765 11747 799
rect 12357 765 12391 799
rect 13001 765 13035 799
rect 13645 765 13679 799
rect 14289 765 14323 799
rect 14933 765 14967 799
rect 15577 765 15611 799
rect 16865 765 16899 799
rect 17509 765 17543 799
rect 18153 765 18187 799
rect 18797 765 18831 799
rect 20085 765 20119 799
<< metal1 >>
rect 552 19066 31372 19088
rect 552 19014 4322 19066
rect 4374 19014 4386 19066
rect 4438 19014 4450 19066
rect 4502 19014 4514 19066
rect 4566 19014 4578 19066
rect 4630 19014 12096 19066
rect 12148 19014 12160 19066
rect 12212 19014 12224 19066
rect 12276 19014 12288 19066
rect 12340 19014 12352 19066
rect 12404 19014 19870 19066
rect 19922 19014 19934 19066
rect 19986 19014 19998 19066
rect 20050 19014 20062 19066
rect 20114 19014 20126 19066
rect 20178 19014 27644 19066
rect 27696 19014 27708 19066
rect 27760 19014 27772 19066
rect 27824 19014 27836 19066
rect 27888 19014 27900 19066
rect 27952 19014 31372 19066
rect 552 18992 31372 19014
rect 14737 18955 14795 18961
rect 14737 18921 14749 18955
rect 14783 18952 14795 18955
rect 14826 18952 14832 18964
rect 14783 18924 14832 18952
rect 14783 18921 14795 18924
rect 14737 18915 14795 18921
rect 14826 18912 14832 18924
rect 14884 18912 14890 18964
rect 16114 18912 16120 18964
rect 16172 18952 16178 18964
rect 17957 18955 18015 18961
rect 17957 18952 17969 18955
rect 16172 18924 17969 18952
rect 16172 18912 16178 18924
rect 17957 18921 17969 18924
rect 18003 18921 18015 18955
rect 17957 18915 18015 18921
rect 10318 18776 10324 18828
rect 10376 18816 10382 18828
rect 10413 18819 10471 18825
rect 10413 18816 10425 18819
rect 10376 18788 10425 18816
rect 10376 18776 10382 18788
rect 10413 18785 10425 18788
rect 10459 18785 10471 18819
rect 10413 18779 10471 18785
rect 11974 18776 11980 18828
rect 12032 18816 12038 18828
rect 12345 18819 12403 18825
rect 12345 18816 12357 18819
rect 12032 18788 12357 18816
rect 12032 18776 12038 18788
rect 12345 18785 12357 18788
rect 12391 18785 12403 18819
rect 12345 18779 12403 18785
rect 12894 18776 12900 18828
rect 12952 18816 12958 18828
rect 12989 18819 13047 18825
rect 12989 18816 13001 18819
rect 12952 18788 13001 18816
rect 12952 18776 12958 18788
rect 12989 18785 13001 18788
rect 13035 18785 13047 18819
rect 12989 18779 13047 18785
rect 13538 18776 13544 18828
rect 13596 18816 13602 18828
rect 13633 18819 13691 18825
rect 13633 18816 13645 18819
rect 13596 18788 13645 18816
rect 13596 18776 13602 18788
rect 13633 18785 13645 18788
rect 13679 18785 13691 18819
rect 13633 18779 13691 18785
rect 14182 18776 14188 18828
rect 14240 18816 14246 18828
rect 14277 18819 14335 18825
rect 14277 18816 14289 18819
rect 14240 18788 14289 18816
rect 14240 18776 14246 18788
rect 14277 18785 14289 18788
rect 14323 18785 14335 18819
rect 14277 18779 14335 18785
rect 14921 18819 14979 18825
rect 14921 18785 14933 18819
rect 14967 18785 14979 18819
rect 14921 18779 14979 18785
rect 17129 18819 17187 18825
rect 17129 18785 17141 18819
rect 17175 18816 17187 18819
rect 17310 18816 17316 18828
rect 17175 18788 17316 18816
rect 17175 18785 17187 18788
rect 17129 18779 17187 18785
rect 14936 18748 14964 18779
rect 17310 18776 17316 18788
rect 17368 18816 17374 18828
rect 17773 18819 17831 18825
rect 17773 18816 17785 18819
rect 17368 18788 17785 18816
rect 17368 18776 17374 18788
rect 17773 18785 17785 18788
rect 17819 18785 17831 18819
rect 17773 18779 17831 18785
rect 18141 18819 18199 18825
rect 18141 18785 18153 18819
rect 18187 18785 18199 18819
rect 18141 18779 18199 18785
rect 15286 18748 15292 18760
rect 14936 18720 15292 18748
rect 15286 18708 15292 18720
rect 15344 18748 15350 18760
rect 15841 18751 15899 18757
rect 15841 18748 15853 18751
rect 15344 18720 15853 18748
rect 15344 18708 15350 18720
rect 15841 18717 15853 18720
rect 15887 18748 15899 18751
rect 16669 18751 16727 18757
rect 16669 18748 16681 18751
rect 15887 18720 16681 18748
rect 15887 18717 15899 18720
rect 15841 18711 15899 18717
rect 16669 18717 16681 18720
rect 16715 18717 16727 18751
rect 16669 18711 16727 18717
rect 17681 18751 17739 18757
rect 17681 18717 17693 18751
rect 17727 18748 17739 18751
rect 18156 18748 18184 18779
rect 22554 18776 22560 18828
rect 22612 18816 22618 18828
rect 22649 18819 22707 18825
rect 22649 18816 22661 18819
rect 22612 18788 22661 18816
rect 22612 18776 22618 18788
rect 22649 18785 22661 18788
rect 22695 18785 22707 18819
rect 22649 18779 22707 18785
rect 17727 18720 18184 18748
rect 17727 18717 17739 18720
rect 17681 18711 17739 18717
rect 16758 18640 16764 18692
rect 16816 18680 16822 18692
rect 18693 18683 18751 18689
rect 18693 18680 18705 18683
rect 16816 18652 18705 18680
rect 16816 18640 16822 18652
rect 18693 18649 18705 18652
rect 18739 18649 18751 18683
rect 18693 18643 18751 18649
rect 842 18572 848 18624
rect 900 18572 906 18624
rect 14366 18572 14372 18624
rect 14424 18612 14430 18624
rect 14461 18615 14519 18621
rect 14461 18612 14473 18615
rect 14424 18584 14473 18612
rect 14424 18572 14430 18584
rect 14461 18581 14473 18584
rect 14507 18581 14519 18615
rect 14461 18575 14519 18581
rect 15194 18572 15200 18624
rect 15252 18572 15258 18624
rect 15378 18572 15384 18624
rect 15436 18612 15442 18624
rect 16117 18615 16175 18621
rect 16117 18612 16129 18615
rect 15436 18584 16129 18612
rect 15436 18572 15442 18584
rect 16117 18581 16129 18584
rect 16163 18581 16175 18615
rect 16117 18575 16175 18581
rect 18230 18572 18236 18624
rect 18288 18572 18294 18624
rect 552 18522 31372 18544
rect 552 18470 3662 18522
rect 3714 18470 3726 18522
rect 3778 18470 3790 18522
rect 3842 18470 3854 18522
rect 3906 18470 3918 18522
rect 3970 18470 11436 18522
rect 11488 18470 11500 18522
rect 11552 18470 11564 18522
rect 11616 18470 11628 18522
rect 11680 18470 11692 18522
rect 11744 18470 19210 18522
rect 19262 18470 19274 18522
rect 19326 18470 19338 18522
rect 19390 18470 19402 18522
rect 19454 18470 19466 18522
rect 19518 18470 26984 18522
rect 27036 18470 27048 18522
rect 27100 18470 27112 18522
rect 27164 18470 27176 18522
rect 27228 18470 27240 18522
rect 27292 18470 31372 18522
rect 552 18448 31372 18470
rect 15286 18368 15292 18420
rect 15344 18368 15350 18420
rect 17310 18417 17316 18420
rect 17267 18411 17316 18417
rect 17267 18408 17279 18411
rect 17223 18380 17279 18408
rect 17267 18377 17279 18380
rect 17313 18377 17316 18411
rect 17267 18371 17316 18377
rect 17310 18368 17316 18371
rect 17368 18408 17374 18420
rect 17405 18411 17463 18417
rect 17405 18408 17417 18411
rect 17368 18380 17417 18408
rect 17368 18368 17374 18380
rect 17405 18377 17417 18380
rect 17451 18377 17463 18411
rect 17405 18371 17463 18377
rect 17494 18368 17500 18420
rect 17552 18408 17558 18420
rect 18049 18411 18107 18417
rect 18049 18408 18061 18411
rect 17552 18380 18061 18408
rect 17552 18368 17558 18380
rect 18049 18377 18061 18380
rect 18095 18377 18107 18411
rect 18049 18371 18107 18377
rect 13817 18275 13875 18281
rect 13817 18241 13829 18275
rect 13863 18272 13875 18275
rect 14182 18272 14188 18284
rect 13863 18244 14188 18272
rect 13863 18241 13875 18244
rect 13817 18235 13875 18241
rect 14182 18232 14188 18244
rect 14240 18232 14246 18284
rect 15473 18275 15531 18281
rect 15473 18241 15485 18275
rect 15519 18272 15531 18275
rect 16390 18272 16396 18284
rect 15519 18244 16396 18272
rect 15519 18241 15531 18244
rect 15473 18235 15531 18241
rect 16390 18232 16396 18244
rect 16448 18232 16454 18284
rect 17126 18232 17132 18284
rect 17184 18272 17190 18284
rect 17497 18275 17555 18281
rect 17497 18272 17509 18275
rect 17184 18244 17509 18272
rect 17184 18232 17190 18244
rect 17497 18241 17509 18244
rect 17543 18241 17555 18275
rect 17497 18235 17555 18241
rect 12710 18164 12716 18216
rect 12768 18204 12774 18216
rect 13541 18207 13599 18213
rect 13541 18204 13553 18207
rect 12768 18176 13553 18204
rect 12768 18164 12774 18176
rect 13541 18173 13553 18176
rect 13587 18173 13599 18207
rect 13541 18167 13599 18173
rect 15838 18164 15844 18216
rect 15896 18164 15902 18216
rect 16758 18164 16764 18216
rect 16816 18204 16822 18216
rect 17405 18207 17463 18213
rect 17405 18204 17417 18207
rect 16816 18176 17417 18204
rect 16816 18164 16822 18176
rect 17405 18173 17417 18176
rect 17451 18204 17463 18207
rect 17865 18207 17923 18213
rect 17865 18204 17877 18207
rect 17451 18176 17877 18204
rect 17451 18173 17463 18176
rect 17405 18167 17463 18173
rect 17865 18173 17877 18176
rect 17911 18173 17923 18207
rect 17865 18167 17923 18173
rect 13648 18108 14306 18136
rect 16882 18108 17356 18136
rect 13648 18080 13676 18108
rect 13630 18028 13636 18080
rect 13688 18028 13694 18080
rect 17328 18068 17356 18108
rect 17678 18068 17684 18080
rect 17328 18040 17684 18068
rect 17678 18028 17684 18040
rect 17736 18028 17742 18080
rect 17770 18028 17776 18080
rect 17828 18028 17834 18080
rect 552 17978 31372 18000
rect 552 17926 4322 17978
rect 4374 17926 4386 17978
rect 4438 17926 4450 17978
rect 4502 17926 4514 17978
rect 4566 17926 4578 17978
rect 4630 17926 12096 17978
rect 12148 17926 12160 17978
rect 12212 17926 12224 17978
rect 12276 17926 12288 17978
rect 12340 17926 12352 17978
rect 12404 17926 19870 17978
rect 19922 17926 19934 17978
rect 19986 17926 19998 17978
rect 20050 17926 20062 17978
rect 20114 17926 20126 17978
rect 20178 17926 27644 17978
rect 27696 17926 27708 17978
rect 27760 17926 27772 17978
rect 27824 17926 27836 17978
rect 27888 17926 27900 17978
rect 27952 17926 31372 17978
rect 552 17904 31372 17926
rect 14108 17836 15332 17864
rect 14108 17805 14136 17836
rect 14093 17799 14151 17805
rect 14093 17765 14105 17799
rect 14139 17765 14151 17799
rect 14734 17796 14740 17808
rect 14093 17759 14151 17765
rect 14476 17768 14740 17796
rect 13630 17688 13636 17740
rect 13688 17688 13694 17740
rect 14476 17737 14504 17768
rect 14734 17756 14740 17768
rect 14792 17756 14798 17808
rect 14921 17799 14979 17805
rect 14921 17765 14933 17799
rect 14967 17796 14979 17799
rect 15194 17796 15200 17808
rect 14967 17768 15200 17796
rect 14967 17765 14979 17768
rect 14921 17759 14979 17765
rect 15194 17756 15200 17768
rect 15252 17756 15258 17808
rect 15304 17796 15332 17836
rect 15838 17824 15844 17876
rect 15896 17864 15902 17876
rect 16117 17867 16175 17873
rect 16117 17864 16129 17867
rect 15896 17836 16129 17864
rect 15896 17824 15902 17836
rect 16117 17833 16129 17836
rect 16163 17833 16175 17867
rect 18230 17864 18236 17876
rect 16117 17827 16175 17833
rect 16224 17836 18236 17864
rect 16224 17796 16252 17836
rect 18230 17824 18236 17836
rect 18288 17824 18294 17876
rect 15304 17768 16252 17796
rect 16577 17799 16635 17805
rect 16577 17765 16589 17799
rect 16623 17796 16635 17799
rect 16623 17768 16988 17796
rect 16623 17765 16635 17768
rect 16577 17759 16635 17765
rect 14461 17731 14519 17737
rect 14461 17697 14473 17731
rect 14507 17697 14519 17731
rect 14461 17691 14519 17697
rect 14642 17688 14648 17740
rect 14700 17688 14706 17740
rect 14829 17731 14887 17737
rect 14829 17697 14841 17731
rect 14875 17728 14887 17731
rect 14875 17700 14964 17728
rect 14875 17697 14887 17700
rect 14829 17691 14887 17697
rect 12253 17663 12311 17669
rect 12253 17629 12265 17663
rect 12299 17629 12311 17663
rect 12253 17623 12311 17629
rect 12268 17524 12296 17623
rect 12526 17620 12532 17672
rect 12584 17620 12590 17672
rect 14277 17663 14335 17669
rect 14277 17629 14289 17663
rect 14323 17629 14335 17663
rect 14277 17623 14335 17629
rect 14292 17592 14320 17623
rect 14366 17620 14372 17672
rect 14424 17620 14430 17672
rect 14642 17592 14648 17604
rect 14292 17564 14648 17592
rect 14642 17552 14648 17564
rect 14700 17552 14706 17604
rect 12710 17524 12716 17536
rect 12268 17496 12716 17524
rect 12710 17484 12716 17496
rect 12768 17484 12774 17536
rect 13998 17484 14004 17536
rect 14056 17484 14062 17536
rect 14182 17484 14188 17536
rect 14240 17524 14246 17536
rect 14277 17527 14335 17533
rect 14277 17524 14289 17527
rect 14240 17496 14289 17524
rect 14240 17484 14246 17496
rect 14277 17493 14289 17496
rect 14323 17493 14335 17527
rect 14936 17524 14964 17700
rect 15010 17688 15016 17740
rect 15068 17688 15074 17740
rect 16485 17731 16543 17737
rect 16485 17697 16497 17731
rect 16531 17728 16543 17731
rect 16850 17728 16856 17740
rect 16531 17700 16856 17728
rect 16531 17697 16543 17700
rect 16485 17691 16543 17697
rect 16850 17688 16856 17700
rect 16908 17688 16914 17740
rect 15286 17620 15292 17672
rect 15344 17620 15350 17672
rect 15841 17663 15899 17669
rect 15841 17629 15853 17663
rect 15887 17629 15899 17663
rect 15841 17623 15899 17629
rect 15197 17595 15255 17601
rect 15197 17561 15209 17595
rect 15243 17592 15255 17595
rect 15856 17592 15884 17623
rect 16298 17620 16304 17672
rect 16356 17660 16362 17672
rect 16960 17669 16988 17768
rect 17954 17756 17960 17808
rect 18012 17756 18018 17808
rect 19058 17756 19064 17808
rect 19116 17796 19122 17808
rect 19116 17768 19288 17796
rect 19116 17756 19122 17768
rect 17126 17688 17132 17740
rect 17184 17728 17190 17740
rect 19260 17737 19288 17768
rect 17221 17731 17279 17737
rect 17221 17728 17233 17731
rect 17184 17700 17233 17728
rect 17184 17688 17190 17700
rect 17221 17697 17233 17700
rect 17267 17728 17279 17731
rect 19245 17731 19303 17737
rect 17267 17700 17448 17728
rect 17267 17697 17279 17700
rect 17221 17691 17279 17697
rect 16669 17663 16727 17669
rect 16669 17660 16681 17663
rect 16356 17632 16681 17660
rect 16356 17620 16362 17632
rect 16669 17629 16681 17632
rect 16715 17629 16727 17663
rect 16669 17623 16727 17629
rect 16945 17663 17003 17669
rect 16945 17629 16957 17663
rect 16991 17660 17003 17663
rect 17310 17660 17316 17672
rect 16991 17632 17316 17660
rect 16991 17629 17003 17632
rect 16945 17623 17003 17629
rect 17310 17620 17316 17632
rect 17368 17620 17374 17672
rect 15243 17564 15884 17592
rect 17420 17592 17448 17700
rect 19245 17697 19257 17731
rect 19291 17697 19303 17731
rect 19245 17691 19303 17697
rect 17586 17620 17592 17672
rect 17644 17660 17650 17672
rect 18969 17663 19027 17669
rect 18969 17660 18981 17663
rect 17644 17632 18981 17660
rect 17644 17620 17650 17632
rect 18969 17629 18981 17632
rect 19015 17629 19027 17663
rect 18969 17623 19027 17629
rect 17497 17595 17555 17601
rect 17497 17592 17509 17595
rect 17420 17564 17509 17592
rect 15243 17561 15255 17564
rect 15197 17555 15255 17561
rect 17497 17561 17509 17564
rect 17543 17561 17555 17595
rect 17497 17555 17555 17561
rect 16758 17524 16764 17536
rect 14936 17496 16764 17524
rect 14277 17487 14335 17493
rect 16758 17484 16764 17496
rect 16816 17524 16822 17536
rect 17037 17527 17095 17533
rect 17037 17524 17049 17527
rect 16816 17496 17049 17524
rect 16816 17484 16822 17496
rect 17037 17493 17049 17496
rect 17083 17493 17095 17527
rect 17037 17487 17095 17493
rect 17402 17484 17408 17536
rect 17460 17484 17466 17536
rect 552 17434 31372 17456
rect 552 17382 3662 17434
rect 3714 17382 3726 17434
rect 3778 17382 3790 17434
rect 3842 17382 3854 17434
rect 3906 17382 3918 17434
rect 3970 17382 11436 17434
rect 11488 17382 11500 17434
rect 11552 17382 11564 17434
rect 11616 17382 11628 17434
rect 11680 17382 11692 17434
rect 11744 17382 19210 17434
rect 19262 17382 19274 17434
rect 19326 17382 19338 17434
rect 19390 17382 19402 17434
rect 19454 17382 19466 17434
rect 19518 17382 26984 17434
rect 27036 17382 27048 17434
rect 27100 17382 27112 17434
rect 27164 17382 27176 17434
rect 27228 17382 27240 17434
rect 27292 17382 31372 17434
rect 552 17360 31372 17382
rect 14642 17280 14648 17332
rect 14700 17320 14706 17332
rect 15102 17320 15108 17332
rect 14700 17292 15108 17320
rect 14700 17280 14706 17292
rect 15102 17280 15108 17292
rect 15160 17320 15166 17332
rect 16298 17320 16304 17332
rect 15160 17292 16304 17320
rect 15160 17280 15166 17292
rect 16298 17280 16304 17292
rect 16356 17280 16362 17332
rect 16758 17280 16764 17332
rect 16816 17280 16822 17332
rect 16850 17280 16856 17332
rect 16908 17280 16914 17332
rect 17586 17280 17592 17332
rect 17644 17280 17650 17332
rect 17770 17280 17776 17332
rect 17828 17280 17834 17332
rect 12710 17212 12716 17264
rect 12768 17252 12774 17264
rect 12768 17224 15056 17252
rect 12768 17212 12774 17224
rect 13630 17144 13636 17196
rect 13688 17184 13694 17196
rect 15028 17193 15056 17224
rect 15013 17187 15071 17193
rect 13688 17156 14872 17184
rect 13688 17144 13694 17156
rect 13722 17076 13728 17128
rect 13780 17076 13786 17128
rect 13998 17076 14004 17128
rect 14056 17076 14062 17128
rect 12710 17008 12716 17060
rect 12768 17048 12774 17060
rect 12805 17051 12863 17057
rect 12805 17048 12817 17051
rect 12768 17020 12817 17048
rect 12768 17008 12774 17020
rect 12805 17017 12817 17020
rect 12851 17017 12863 17051
rect 14844 17048 14872 17156
rect 15013 17153 15025 17187
rect 15059 17153 15071 17187
rect 15013 17147 15071 17153
rect 15286 17144 15292 17196
rect 15344 17144 15350 17196
rect 16776 17184 16804 17280
rect 17405 17187 17463 17193
rect 17405 17184 17417 17187
rect 16776 17156 17417 17184
rect 17405 17153 17417 17156
rect 17451 17153 17463 17187
rect 17405 17147 17463 17153
rect 18322 17144 18328 17196
rect 18380 17144 18386 17196
rect 14921 17119 14979 17125
rect 14921 17085 14933 17119
rect 14967 17116 14979 17119
rect 17954 17116 17960 17128
rect 14967 17088 15056 17116
rect 14967 17085 14979 17088
rect 14921 17079 14979 17085
rect 15028 17048 15056 17088
rect 17328 17088 17960 17116
rect 17328 17060 17356 17088
rect 17954 17076 17960 17088
rect 18012 17076 18018 17128
rect 18141 17119 18199 17125
rect 18141 17085 18153 17119
rect 18187 17116 18199 17119
rect 18340 17116 18368 17144
rect 18509 17119 18567 17125
rect 18509 17116 18521 17119
rect 18187 17088 18521 17116
rect 18187 17085 18199 17088
rect 18141 17079 18199 17085
rect 18509 17085 18521 17088
rect 18555 17085 18567 17119
rect 18509 17079 18567 17085
rect 15378 17048 15384 17060
rect 14844 17020 14964 17048
rect 15028 17020 15384 17048
rect 12805 17011 12863 17017
rect 13814 16940 13820 16992
rect 13872 16940 13878 16992
rect 14182 16940 14188 16992
rect 14240 16940 14246 16992
rect 14826 16940 14832 16992
rect 14884 16940 14890 16992
rect 14936 16980 14964 17020
rect 15378 17008 15384 17020
rect 15436 17008 15442 17060
rect 17310 17048 17316 17060
rect 15672 17020 15778 17048
rect 16592 17020 17316 17048
rect 15672 16980 15700 17020
rect 16592 16980 16620 17020
rect 17310 17008 17316 17020
rect 17368 17008 17374 17060
rect 17402 17008 17408 17060
rect 17460 17048 17466 17060
rect 17678 17048 17684 17060
rect 17460 17020 17684 17048
rect 17460 17008 17466 17020
rect 17678 17008 17684 17020
rect 17736 17048 17742 17060
rect 18325 17051 18383 17057
rect 18325 17048 18337 17051
rect 17736 17020 18337 17048
rect 17736 17008 17742 17020
rect 18325 17017 18337 17020
rect 18371 17017 18383 17051
rect 18325 17011 18383 17017
rect 14936 16952 16620 16980
rect 16666 16940 16672 16992
rect 16724 16980 16730 16992
rect 17494 16980 17500 16992
rect 16724 16952 17500 16980
rect 16724 16940 16730 16952
rect 17494 16940 17500 16952
rect 17552 16980 17558 16992
rect 17773 16983 17831 16989
rect 17773 16980 17785 16983
rect 17552 16952 17785 16980
rect 17552 16940 17558 16952
rect 17773 16949 17785 16952
rect 17819 16949 17831 16983
rect 17773 16943 17831 16949
rect 552 16890 31372 16912
rect 552 16838 4322 16890
rect 4374 16838 4386 16890
rect 4438 16838 4450 16890
rect 4502 16838 4514 16890
rect 4566 16838 4578 16890
rect 4630 16838 12096 16890
rect 12148 16838 12160 16890
rect 12212 16838 12224 16890
rect 12276 16838 12288 16890
rect 12340 16838 12352 16890
rect 12404 16838 19870 16890
rect 19922 16838 19934 16890
rect 19986 16838 19998 16890
rect 20050 16838 20062 16890
rect 20114 16838 20126 16890
rect 20178 16838 27644 16890
rect 27696 16838 27708 16890
rect 27760 16838 27772 16890
rect 27824 16838 27836 16890
rect 27888 16838 27900 16890
rect 27952 16838 31372 16890
rect 552 16816 31372 16838
rect 14182 16736 14188 16788
rect 14240 16776 14246 16788
rect 15013 16779 15071 16785
rect 15013 16776 15025 16779
rect 14240 16748 15025 16776
rect 14240 16736 14246 16748
rect 15013 16745 15025 16748
rect 15059 16745 15071 16779
rect 15013 16739 15071 16745
rect 15470 16736 15476 16788
rect 15528 16776 15534 16788
rect 15528 16748 19288 16776
rect 15528 16736 15534 16748
rect 14461 16711 14519 16717
rect 14461 16677 14473 16711
rect 14507 16708 14519 16711
rect 15488 16708 15516 16736
rect 14507 16680 15516 16708
rect 16209 16711 16267 16717
rect 14507 16677 14519 16680
rect 14461 16671 14519 16677
rect 16209 16677 16221 16711
rect 16255 16708 16267 16711
rect 16666 16708 16672 16720
rect 16255 16680 16672 16708
rect 16255 16677 16267 16680
rect 16209 16671 16267 16677
rect 16666 16668 16672 16680
rect 16724 16668 16730 16720
rect 17126 16708 17132 16720
rect 16868 16680 17132 16708
rect 12526 16600 12532 16652
rect 12584 16640 12590 16652
rect 14553 16643 14611 16649
rect 14553 16640 14565 16643
rect 12584 16612 14565 16640
rect 12584 16600 12590 16612
rect 14553 16609 14565 16612
rect 14599 16609 14611 16643
rect 14553 16603 14611 16609
rect 14826 16600 14832 16652
rect 14884 16600 14890 16652
rect 14921 16643 14979 16649
rect 14921 16609 14933 16643
rect 14967 16640 14979 16643
rect 15194 16640 15200 16652
rect 14967 16612 15200 16640
rect 14967 16609 14979 16612
rect 14921 16603 14979 16609
rect 15194 16600 15200 16612
rect 15252 16600 15258 16652
rect 15289 16643 15347 16649
rect 15289 16609 15301 16643
rect 15335 16640 15347 16643
rect 15473 16643 15531 16649
rect 15473 16640 15485 16643
rect 15335 16612 15485 16640
rect 15335 16609 15347 16612
rect 15289 16603 15347 16609
rect 15473 16609 15485 16612
rect 15519 16609 15531 16643
rect 15473 16603 15531 16609
rect 15562 16600 15568 16652
rect 15620 16600 15626 16652
rect 16485 16643 16543 16649
rect 16485 16640 16497 16643
rect 15672 16612 16497 16640
rect 12710 16532 12716 16584
rect 12768 16532 12774 16584
rect 14844 16572 14872 16600
rect 15672 16572 15700 16612
rect 16485 16609 16497 16612
rect 16531 16609 16543 16643
rect 16485 16603 16543 16609
rect 16574 16600 16580 16652
rect 16632 16640 16638 16652
rect 16868 16649 16896 16680
rect 17126 16668 17132 16680
rect 17184 16668 17190 16720
rect 17310 16668 17316 16720
rect 17368 16708 17374 16720
rect 19260 16717 19288 16748
rect 19245 16711 19303 16717
rect 17368 16680 17710 16708
rect 17368 16668 17374 16680
rect 19245 16677 19257 16711
rect 19291 16677 19303 16711
rect 19245 16671 19303 16677
rect 16853 16643 16911 16649
rect 16853 16640 16865 16643
rect 16632 16612 16865 16640
rect 16632 16600 16638 16612
rect 16853 16609 16865 16612
rect 16899 16609 16911 16643
rect 16853 16603 16911 16609
rect 17034 16600 17040 16652
rect 17092 16600 17098 16652
rect 17218 16600 17224 16652
rect 17276 16600 17282 16652
rect 19150 16600 19156 16652
rect 19208 16600 19214 16652
rect 14844 16544 15700 16572
rect 17236 16572 17264 16600
rect 17405 16575 17463 16581
rect 17405 16572 17417 16575
rect 17236 16544 17417 16572
rect 17405 16541 17417 16544
rect 17451 16541 17463 16575
rect 17405 16535 17463 16541
rect 18874 16532 18880 16584
rect 18932 16532 18938 16584
rect 13998 16464 14004 16516
rect 14056 16504 14062 16516
rect 15562 16504 15568 16516
rect 14056 16476 15568 16504
rect 14056 16464 14062 16476
rect 15562 16464 15568 16476
rect 15620 16464 15626 16516
rect 16577 16507 16635 16513
rect 16577 16473 16589 16507
rect 16623 16504 16635 16507
rect 16942 16504 16948 16516
rect 16623 16476 16948 16504
rect 16623 16473 16635 16476
rect 16577 16467 16635 16473
rect 16942 16464 16948 16476
rect 17000 16504 17006 16516
rect 17129 16507 17187 16513
rect 17129 16504 17141 16507
rect 17000 16476 17141 16504
rect 17000 16464 17006 16476
rect 17129 16473 17141 16476
rect 17175 16473 17187 16507
rect 17129 16467 17187 16473
rect 19150 16464 19156 16516
rect 19208 16504 19214 16516
rect 20533 16507 20591 16513
rect 20533 16504 20545 16507
rect 19208 16476 20545 16504
rect 19208 16464 19214 16476
rect 20533 16473 20545 16476
rect 20579 16473 20591 16507
rect 20533 16467 20591 16473
rect 15197 16439 15255 16445
rect 15197 16405 15209 16439
rect 15243 16436 15255 16439
rect 15838 16436 15844 16448
rect 15243 16408 15844 16436
rect 15243 16405 15255 16408
rect 15197 16399 15255 16405
rect 15838 16396 15844 16408
rect 15896 16396 15902 16448
rect 16666 16396 16672 16448
rect 16724 16396 16730 16448
rect 16761 16439 16819 16445
rect 16761 16405 16773 16439
rect 16807 16436 16819 16439
rect 17034 16436 17040 16448
rect 16807 16408 17040 16436
rect 16807 16405 16819 16408
rect 16761 16399 16819 16405
rect 17034 16396 17040 16408
rect 17092 16396 17098 16448
rect 552 16346 31372 16368
rect 552 16294 3662 16346
rect 3714 16294 3726 16346
rect 3778 16294 3790 16346
rect 3842 16294 3854 16346
rect 3906 16294 3918 16346
rect 3970 16294 11436 16346
rect 11488 16294 11500 16346
rect 11552 16294 11564 16346
rect 11616 16294 11628 16346
rect 11680 16294 11692 16346
rect 11744 16294 19210 16346
rect 19262 16294 19274 16346
rect 19326 16294 19338 16346
rect 19390 16294 19402 16346
rect 19454 16294 19466 16346
rect 19518 16294 26984 16346
rect 27036 16294 27048 16346
rect 27100 16294 27112 16346
rect 27164 16294 27176 16346
rect 27228 16294 27240 16346
rect 27292 16294 31372 16346
rect 552 16272 31372 16294
rect 12802 16192 12808 16244
rect 12860 16232 12866 16244
rect 12897 16235 12955 16241
rect 12897 16232 12909 16235
rect 12860 16204 12909 16232
rect 12860 16192 12866 16204
rect 12897 16201 12909 16204
rect 12943 16232 12955 16235
rect 14550 16232 14556 16244
rect 12943 16204 14556 16232
rect 12943 16201 12955 16204
rect 12897 16195 12955 16201
rect 14550 16192 14556 16204
rect 14608 16192 14614 16244
rect 15470 16192 15476 16244
rect 15528 16192 15534 16244
rect 18325 16235 18383 16241
rect 18325 16201 18337 16235
rect 18371 16232 18383 16235
rect 19334 16232 19340 16244
rect 18371 16204 19340 16232
rect 18371 16201 18383 16204
rect 18325 16195 18383 16201
rect 13998 16124 14004 16176
rect 14056 16124 14062 16176
rect 18230 16164 18236 16176
rect 16868 16136 18236 16164
rect 13909 16099 13967 16105
rect 13909 16065 13921 16099
rect 13955 16096 13967 16099
rect 14016 16096 14044 16124
rect 13955 16068 14044 16096
rect 13955 16065 13967 16068
rect 13909 16059 13967 16065
rect 14366 16056 14372 16108
rect 14424 16096 14430 16108
rect 15746 16096 15752 16108
rect 14424 16068 15752 16096
rect 14424 16056 14430 16068
rect 15746 16056 15752 16068
rect 15804 16096 15810 16108
rect 16868 16096 16896 16136
rect 18230 16124 18236 16136
rect 18288 16124 18294 16176
rect 18340 16096 18368 16195
rect 19334 16192 19340 16204
rect 19392 16192 19398 16244
rect 15804 16068 16896 16096
rect 15804 16056 15810 16068
rect 12986 15988 12992 16040
rect 13044 16028 13050 16040
rect 13265 16031 13323 16037
rect 13265 16028 13277 16031
rect 13044 16000 13277 16028
rect 13044 15988 13050 16000
rect 13265 15997 13277 16000
rect 13311 15997 13323 16031
rect 13265 15991 13323 15997
rect 13722 15988 13728 16040
rect 13780 15988 13786 16040
rect 13814 15988 13820 16040
rect 13872 15988 13878 16040
rect 13998 15988 14004 16040
rect 14056 15988 14062 16040
rect 16868 16037 16896 16068
rect 17144 16068 18368 16096
rect 16853 16031 16911 16037
rect 16853 15997 16865 16031
rect 16899 15997 16911 16031
rect 16853 15991 16911 15997
rect 17034 15988 17040 16040
rect 17092 16028 17098 16040
rect 17144 16037 17172 16068
rect 17129 16031 17187 16037
rect 17129 16028 17141 16031
rect 17092 16000 17141 16028
rect 17092 15988 17098 16000
rect 17129 15997 17141 16000
rect 17175 15997 17187 16031
rect 17129 15991 17187 15997
rect 17218 15988 17224 16040
rect 17276 16028 17282 16040
rect 17957 16031 18015 16037
rect 17957 16028 17969 16031
rect 17276 16000 17969 16028
rect 17276 15988 17282 16000
rect 17957 15997 17969 16000
rect 18003 15997 18015 16031
rect 17957 15991 18015 15997
rect 13832 15960 13860 15988
rect 14366 15960 14372 15972
rect 13832 15932 14372 15960
rect 14366 15920 14372 15932
rect 14424 15920 14430 15972
rect 16758 15920 16764 15972
rect 16816 15920 16822 15972
rect 16945 15963 17003 15969
rect 16945 15929 16957 15963
rect 16991 15960 17003 15963
rect 18046 15960 18052 15972
rect 16991 15932 18052 15960
rect 16991 15929 17003 15932
rect 16945 15923 17003 15929
rect 17144 15904 17172 15932
rect 18046 15920 18052 15932
rect 18104 15960 18110 15972
rect 18322 15969 18328 15972
rect 18309 15963 18328 15969
rect 18104 15932 18276 15960
rect 18104 15920 18110 15932
rect 12526 15852 12532 15904
rect 12584 15892 12590 15904
rect 12713 15895 12771 15901
rect 12713 15892 12725 15895
rect 12584 15864 12725 15892
rect 12584 15852 12590 15864
rect 12713 15861 12725 15864
rect 12759 15861 12771 15895
rect 12713 15855 12771 15861
rect 12897 15895 12955 15901
rect 12897 15861 12909 15895
rect 12943 15892 12955 15895
rect 13541 15895 13599 15901
rect 13541 15892 13553 15895
rect 12943 15864 13553 15892
rect 12943 15861 12955 15864
rect 12897 15855 12955 15861
rect 13541 15861 13553 15864
rect 13587 15861 13599 15895
rect 13541 15855 13599 15861
rect 16850 15852 16856 15904
rect 16908 15892 16914 15904
rect 17126 15892 17132 15904
rect 16908 15864 17132 15892
rect 16908 15852 16914 15864
rect 17126 15852 17132 15864
rect 17184 15852 17190 15904
rect 17310 15852 17316 15904
rect 17368 15852 17374 15904
rect 17402 15852 17408 15904
rect 17460 15852 17466 15904
rect 17586 15852 17592 15904
rect 17644 15892 17650 15904
rect 18141 15895 18199 15901
rect 18141 15892 18153 15895
rect 17644 15864 18153 15892
rect 17644 15852 17650 15864
rect 18141 15861 18153 15864
rect 18187 15861 18199 15895
rect 18248 15892 18276 15932
rect 18309 15929 18321 15963
rect 18309 15923 18328 15929
rect 18322 15920 18328 15923
rect 18380 15920 18386 15972
rect 18509 15963 18567 15969
rect 18509 15929 18521 15963
rect 18555 15929 18567 15963
rect 18509 15923 18567 15929
rect 18524 15892 18552 15923
rect 18248 15864 18552 15892
rect 18141 15855 18199 15861
rect 552 15802 31372 15824
rect 552 15750 4322 15802
rect 4374 15750 4386 15802
rect 4438 15750 4450 15802
rect 4502 15750 4514 15802
rect 4566 15750 4578 15802
rect 4630 15750 12096 15802
rect 12148 15750 12160 15802
rect 12212 15750 12224 15802
rect 12276 15750 12288 15802
rect 12340 15750 12352 15802
rect 12404 15750 19870 15802
rect 19922 15750 19934 15802
rect 19986 15750 19998 15802
rect 20050 15750 20062 15802
rect 20114 15750 20126 15802
rect 20178 15750 27644 15802
rect 27696 15750 27708 15802
rect 27760 15750 27772 15802
rect 27824 15750 27836 15802
rect 27888 15750 27900 15802
rect 27952 15750 31372 15802
rect 552 15728 31372 15750
rect 13998 15648 14004 15700
rect 14056 15648 14062 15700
rect 14090 15648 14096 15700
rect 14148 15688 14154 15700
rect 14461 15691 14519 15697
rect 14461 15688 14473 15691
rect 14148 15660 14473 15688
rect 14148 15648 14154 15660
rect 14461 15657 14473 15660
rect 14507 15688 14519 15691
rect 14734 15688 14740 15700
rect 14507 15660 14740 15688
rect 14507 15657 14519 15660
rect 14461 15651 14519 15657
rect 14734 15648 14740 15660
rect 14792 15648 14798 15700
rect 15197 15691 15255 15697
rect 15197 15657 15209 15691
rect 15243 15688 15255 15691
rect 16942 15688 16948 15700
rect 15243 15660 16620 15688
rect 15243 15657 15255 15660
rect 15197 15651 15255 15657
rect 12526 15580 12532 15632
rect 12584 15580 12590 15632
rect 14016 15620 14044 15648
rect 14645 15623 14703 15629
rect 14645 15620 14657 15623
rect 14016 15592 14657 15620
rect 14645 15589 14657 15592
rect 14691 15620 14703 15623
rect 14691 15592 15056 15620
rect 14691 15589 14703 15592
rect 14645 15583 14703 15589
rect 13630 15512 13636 15564
rect 13688 15512 13694 15564
rect 13814 15512 13820 15564
rect 13872 15552 13878 15564
rect 14277 15555 14335 15561
rect 14277 15552 14289 15555
rect 13872 15524 14289 15552
rect 13872 15512 13878 15524
rect 14277 15521 14289 15524
rect 14323 15521 14335 15555
rect 14277 15515 14335 15521
rect 12253 15487 12311 15493
rect 12253 15453 12265 15487
rect 12299 15453 12311 15487
rect 12253 15447 12311 15453
rect 12268 15348 12296 15447
rect 12986 15444 12992 15496
rect 13044 15484 13050 15496
rect 14093 15487 14151 15493
rect 14093 15484 14105 15487
rect 13044 15456 14105 15484
rect 13044 15444 13050 15456
rect 14093 15453 14105 15456
rect 14139 15453 14151 15487
rect 14292 15484 14320 15515
rect 14366 15512 14372 15564
rect 14424 15512 14430 15564
rect 14458 15512 14464 15564
rect 14516 15552 14522 15564
rect 14737 15555 14795 15561
rect 14660 15552 14749 15555
rect 14516 15527 14749 15552
rect 14516 15524 14688 15527
rect 14516 15512 14522 15524
rect 14737 15521 14749 15527
rect 14783 15521 14795 15555
rect 14737 15515 14795 15521
rect 14918 15512 14924 15564
rect 14976 15512 14982 15564
rect 15028 15561 15056 15592
rect 15838 15580 15844 15632
rect 15896 15580 15902 15632
rect 15013 15555 15071 15561
rect 15013 15521 15025 15555
rect 15059 15552 15071 15555
rect 15470 15552 15476 15564
rect 15059 15524 15476 15552
rect 15059 15521 15071 15524
rect 15013 15515 15071 15521
rect 15470 15512 15476 15524
rect 15528 15512 15534 15564
rect 15746 15512 15752 15564
rect 15804 15512 15810 15564
rect 15562 15484 15568 15496
rect 14292 15456 15568 15484
rect 14093 15447 14151 15453
rect 15562 15444 15568 15456
rect 15620 15444 15626 15496
rect 15856 15484 15884 15580
rect 15930 15512 15936 15564
rect 15988 15512 15994 15564
rect 16482 15512 16488 15564
rect 16540 15512 16546 15564
rect 16592 15561 16620 15660
rect 16776 15660 16948 15688
rect 16776 15629 16804 15660
rect 16942 15648 16948 15660
rect 17000 15648 17006 15700
rect 17494 15648 17500 15700
rect 17552 15648 17558 15700
rect 18874 15688 18880 15700
rect 17880 15660 18880 15688
rect 16761 15623 16819 15629
rect 16761 15589 16773 15623
rect 16807 15589 16819 15623
rect 17512 15620 17540 15648
rect 17880 15620 17908 15660
rect 18874 15648 18880 15660
rect 18932 15648 18938 15700
rect 19334 15648 19340 15700
rect 19392 15648 19398 15700
rect 16761 15583 16819 15589
rect 16868 15592 17540 15620
rect 17604 15592 17908 15620
rect 16577 15555 16635 15561
rect 16577 15521 16589 15555
rect 16623 15552 16635 15555
rect 16666 15552 16672 15564
rect 16623 15524 16672 15552
rect 16623 15521 16635 15524
rect 16577 15515 16635 15521
rect 16666 15512 16672 15524
rect 16724 15512 16730 15564
rect 16868 15561 16896 15592
rect 16853 15555 16911 15561
rect 16853 15521 16865 15555
rect 16899 15521 16911 15555
rect 16853 15515 16911 15521
rect 17037 15555 17095 15561
rect 17037 15521 17049 15555
rect 17083 15521 17095 15555
rect 17037 15515 17095 15521
rect 17052 15484 17080 15515
rect 17126 15512 17132 15564
rect 17184 15512 17190 15564
rect 17221 15555 17279 15561
rect 17221 15521 17233 15555
rect 17267 15552 17279 15555
rect 17402 15552 17408 15564
rect 17267 15524 17408 15552
rect 17267 15521 17279 15524
rect 17221 15515 17279 15521
rect 17402 15512 17408 15524
rect 17460 15512 17466 15564
rect 17604 15552 17632 15592
rect 17954 15580 17960 15632
rect 18012 15620 18018 15632
rect 18322 15620 18328 15632
rect 18012 15592 18328 15620
rect 18012 15580 18018 15592
rect 18322 15580 18328 15592
rect 18380 15580 18386 15632
rect 17512 15524 17632 15552
rect 17512 15493 17540 15524
rect 15856 15456 17080 15484
rect 17497 15487 17555 15493
rect 17497 15453 17509 15487
rect 17543 15453 17555 15487
rect 17497 15447 17555 15453
rect 17589 15487 17647 15493
rect 17589 15453 17601 15487
rect 17635 15453 17647 15487
rect 17589 15447 17647 15453
rect 13906 15376 13912 15428
rect 13964 15416 13970 15428
rect 14918 15416 14924 15428
rect 13964 15388 14924 15416
rect 13964 15376 13970 15388
rect 14918 15376 14924 15388
rect 14976 15376 14982 15428
rect 15194 15376 15200 15428
rect 15252 15416 15258 15428
rect 16301 15419 16359 15425
rect 16301 15416 16313 15419
rect 15252 15388 16313 15416
rect 15252 15376 15258 15388
rect 16301 15385 16313 15388
rect 16347 15385 16359 15419
rect 16301 15379 16359 15385
rect 16482 15376 16488 15428
rect 16540 15416 16546 15428
rect 16540 15388 17448 15416
rect 16540 15376 16546 15388
rect 12710 15348 12716 15360
rect 12268 15320 12716 15348
rect 12710 15308 12716 15320
rect 12768 15308 12774 15360
rect 14734 15308 14740 15360
rect 14792 15308 14798 15360
rect 16761 15351 16819 15357
rect 16761 15317 16773 15351
rect 16807 15348 16819 15351
rect 17034 15348 17040 15360
rect 16807 15320 17040 15348
rect 16807 15317 16819 15320
rect 16761 15311 16819 15317
rect 17034 15308 17040 15320
rect 17092 15308 17098 15360
rect 17420 15348 17448 15388
rect 17604 15348 17632 15447
rect 17862 15444 17868 15496
rect 17920 15444 17926 15496
rect 19058 15348 19064 15360
rect 17420 15320 19064 15348
rect 19058 15308 19064 15320
rect 19116 15308 19122 15360
rect 552 15258 31372 15280
rect 552 15206 3662 15258
rect 3714 15206 3726 15258
rect 3778 15206 3790 15258
rect 3842 15206 3854 15258
rect 3906 15206 3918 15258
rect 3970 15206 11436 15258
rect 11488 15206 11500 15258
rect 11552 15206 11564 15258
rect 11616 15206 11628 15258
rect 11680 15206 11692 15258
rect 11744 15206 19210 15258
rect 19262 15206 19274 15258
rect 19326 15206 19338 15258
rect 19390 15206 19402 15258
rect 19454 15206 19466 15258
rect 19518 15206 26984 15258
rect 27036 15206 27048 15258
rect 27100 15206 27112 15258
rect 27164 15206 27176 15258
rect 27228 15206 27240 15258
rect 27292 15206 31372 15258
rect 552 15184 31372 15206
rect 12618 15104 12624 15156
rect 12676 15144 12682 15156
rect 12676 15116 13860 15144
rect 12676 15104 12682 15116
rect 13832 15088 13860 15116
rect 14734 15104 14740 15156
rect 14792 15144 14798 15156
rect 15749 15147 15807 15153
rect 15749 15144 15761 15147
rect 14792 15116 15761 15144
rect 14792 15104 14798 15116
rect 15749 15113 15761 15116
rect 15795 15113 15807 15147
rect 15749 15107 15807 15113
rect 15930 15104 15936 15156
rect 15988 15144 15994 15156
rect 16393 15147 16451 15153
rect 16393 15144 16405 15147
rect 15988 15116 16405 15144
rect 15988 15104 15994 15116
rect 16393 15113 16405 15116
rect 16439 15113 16451 15147
rect 16393 15107 16451 15113
rect 16577 15147 16635 15153
rect 16577 15113 16589 15147
rect 16623 15144 16635 15147
rect 17034 15144 17040 15156
rect 16623 15116 17040 15144
rect 16623 15113 16635 15116
rect 16577 15107 16635 15113
rect 17034 15104 17040 15116
rect 17092 15104 17098 15156
rect 17494 15104 17500 15156
rect 17552 15104 17558 15156
rect 17681 15147 17739 15153
rect 17681 15113 17693 15147
rect 17727 15144 17739 15147
rect 17862 15144 17868 15156
rect 17727 15116 17868 15144
rect 17727 15113 17739 15116
rect 17681 15107 17739 15113
rect 17862 15104 17868 15116
rect 17920 15104 17926 15156
rect 12526 15036 12532 15088
rect 12584 15076 12590 15088
rect 13722 15076 13728 15088
rect 12584 15048 13728 15076
rect 12584 15036 12590 15048
rect 13722 15036 13728 15048
rect 13780 15036 13786 15088
rect 13814 15036 13820 15088
rect 13872 15076 13878 15088
rect 14366 15076 14372 15088
rect 13872 15048 14372 15076
rect 13872 15036 13878 15048
rect 14366 15036 14372 15048
rect 14424 15036 14430 15088
rect 15565 15079 15623 15085
rect 15565 15076 15577 15079
rect 15120 15048 15577 15076
rect 15120 15017 15148 15048
rect 15565 15045 15577 15048
rect 15611 15045 15623 15079
rect 15565 15039 15623 15045
rect 17126 15036 17132 15088
rect 17184 15076 17190 15088
rect 17586 15076 17592 15088
rect 17184 15048 17592 15076
rect 17184 15036 17190 15048
rect 17586 15036 17592 15048
rect 17644 15036 17650 15088
rect 15105 15011 15163 15017
rect 15105 15008 15117 15011
rect 12360 14980 15117 15008
rect 12360 14949 12388 14980
rect 12345 14943 12403 14949
rect 12345 14909 12357 14943
rect 12391 14909 12403 14943
rect 12345 14903 12403 14909
rect 12526 14900 12532 14952
rect 12584 14900 12590 14952
rect 12618 14900 12624 14952
rect 12676 14900 12682 14952
rect 12713 14943 12771 14949
rect 12713 14909 12725 14943
rect 12759 14940 12771 14943
rect 12802 14940 12808 14952
rect 12759 14912 12808 14940
rect 12759 14909 12771 14912
rect 12713 14903 12771 14909
rect 12802 14900 12808 14912
rect 12860 14900 12866 14952
rect 12897 14943 12955 14949
rect 12897 14909 12909 14943
rect 12943 14909 12955 14943
rect 12897 14903 12955 14909
rect 12912 14872 12940 14903
rect 12986 14900 12992 14952
rect 13044 14900 13050 14952
rect 13556 14949 13584 14980
rect 15105 14977 15117 14980
rect 15151 14977 15163 15011
rect 15105 14971 15163 14977
rect 15289 15011 15347 15017
rect 15289 14977 15301 15011
rect 15335 15008 15347 15011
rect 15746 15008 15752 15020
rect 15335 14980 15752 15008
rect 15335 14977 15347 14980
rect 15289 14971 15347 14977
rect 15746 14968 15752 14980
rect 15804 14968 15810 15020
rect 13081 14943 13139 14949
rect 13081 14909 13093 14943
rect 13127 14909 13139 14943
rect 13081 14903 13139 14909
rect 13541 14943 13599 14949
rect 13541 14909 13553 14943
rect 13587 14909 13599 14943
rect 13541 14903 13599 14909
rect 13633 14943 13691 14949
rect 13633 14909 13645 14943
rect 13679 14940 13691 14943
rect 13722 14940 13728 14952
rect 13679 14912 13728 14940
rect 13679 14909 13691 14912
rect 13633 14903 13691 14909
rect 12636 14844 12940 14872
rect 13096 14872 13124 14903
rect 13722 14900 13728 14912
rect 13780 14900 13786 14952
rect 13906 14900 13912 14952
rect 13964 14900 13970 14952
rect 14458 14900 14464 14952
rect 14516 14940 14522 14952
rect 14737 14943 14795 14949
rect 14737 14940 14749 14943
rect 14516 14912 14749 14940
rect 14516 14900 14522 14912
rect 14737 14909 14749 14912
rect 14783 14909 14795 14943
rect 14737 14903 14795 14909
rect 14185 14875 14243 14881
rect 14185 14872 14197 14875
rect 13096 14844 14197 14872
rect 12636 14813 12664 14844
rect 14185 14841 14197 14844
rect 14231 14841 14243 14875
rect 14752 14872 14780 14903
rect 15194 14900 15200 14952
rect 15252 14900 15258 14952
rect 15378 14900 15384 14952
rect 15436 14900 15442 14952
rect 15470 14900 15476 14952
rect 15528 14940 15534 14952
rect 16850 14940 16856 14952
rect 15528 14912 15976 14940
rect 15528 14900 15534 14912
rect 15948 14881 15976 14912
rect 16776 14912 16856 14940
rect 16776 14881 16804 14912
rect 16850 14900 16856 14912
rect 16908 14900 16914 14952
rect 17037 14943 17095 14949
rect 17037 14909 17049 14943
rect 17083 14940 17095 14943
rect 17678 14940 17684 14952
rect 17083 14912 17684 14940
rect 17083 14909 17095 14912
rect 17037 14903 17095 14909
rect 17678 14900 17684 14912
rect 17736 14900 17742 14952
rect 15717 14875 15775 14881
rect 15717 14872 15729 14875
rect 14752 14844 15729 14872
rect 14185 14835 14243 14841
rect 15717 14841 15729 14844
rect 15763 14841 15775 14875
rect 15717 14835 15775 14841
rect 15933 14875 15991 14881
rect 15933 14841 15945 14875
rect 15979 14841 15991 14875
rect 15933 14835 15991 14841
rect 16761 14875 16819 14881
rect 16761 14841 16773 14875
rect 16807 14841 16819 14875
rect 17218 14872 17224 14884
rect 16761 14835 16819 14841
rect 16868 14844 17224 14872
rect 12621 14807 12679 14813
rect 12621 14773 12633 14807
rect 12667 14773 12679 14807
rect 12621 14767 12679 14773
rect 12986 14764 12992 14816
rect 13044 14804 13050 14816
rect 13357 14807 13415 14813
rect 13357 14804 13369 14807
rect 13044 14776 13369 14804
rect 13044 14764 13050 14776
rect 13357 14773 13369 14776
rect 13403 14773 13415 14807
rect 13357 14767 13415 14773
rect 13725 14807 13783 14813
rect 13725 14773 13737 14807
rect 13771 14804 13783 14807
rect 13814 14804 13820 14816
rect 13771 14776 13820 14804
rect 13771 14773 13783 14776
rect 13725 14767 13783 14773
rect 13814 14764 13820 14776
rect 13872 14764 13878 14816
rect 13909 14807 13967 14813
rect 13909 14773 13921 14807
rect 13955 14804 13967 14807
rect 13998 14804 14004 14816
rect 13955 14776 14004 14804
rect 13955 14773 13967 14776
rect 13909 14767 13967 14773
rect 13998 14764 14004 14776
rect 14056 14764 14062 14816
rect 14918 14764 14924 14816
rect 14976 14764 14982 14816
rect 15194 14764 15200 14816
rect 15252 14804 15258 14816
rect 15562 14804 15568 14816
rect 15252 14776 15568 14804
rect 15252 14764 15258 14776
rect 15562 14764 15568 14776
rect 15620 14804 15626 14816
rect 15838 14804 15844 14816
rect 15620 14776 15844 14804
rect 15620 14764 15626 14776
rect 15838 14764 15844 14776
rect 15896 14764 15902 14816
rect 16577 14807 16635 14813
rect 16577 14773 16589 14807
rect 16623 14804 16635 14807
rect 16868 14804 16896 14844
rect 17218 14832 17224 14844
rect 17276 14832 17282 14884
rect 17310 14832 17316 14884
rect 17368 14872 17374 14884
rect 17497 14875 17555 14881
rect 17497 14872 17509 14875
rect 17368 14844 17509 14872
rect 17368 14832 17374 14844
rect 17497 14841 17509 14844
rect 17543 14841 17555 14875
rect 17497 14835 17555 14841
rect 16623 14776 16896 14804
rect 16623 14773 16635 14776
rect 16577 14767 16635 14773
rect 16942 14764 16948 14816
rect 17000 14764 17006 14816
rect 552 14714 31372 14736
rect 552 14662 4322 14714
rect 4374 14662 4386 14714
rect 4438 14662 4450 14714
rect 4502 14662 4514 14714
rect 4566 14662 4578 14714
rect 4630 14662 12096 14714
rect 12148 14662 12160 14714
rect 12212 14662 12224 14714
rect 12276 14662 12288 14714
rect 12340 14662 12352 14714
rect 12404 14662 19870 14714
rect 19922 14662 19934 14714
rect 19986 14662 19998 14714
rect 20050 14662 20062 14714
rect 20114 14662 20126 14714
rect 20178 14662 27644 14714
rect 27696 14662 27708 14714
rect 27760 14662 27772 14714
rect 27824 14662 27836 14714
rect 27888 14662 27900 14714
rect 27952 14662 31372 14714
rect 552 14640 31372 14662
rect 14458 14560 14464 14612
rect 14516 14560 14522 14612
rect 14763 14603 14821 14609
rect 14763 14569 14775 14603
rect 14809 14600 14821 14603
rect 14918 14600 14924 14612
rect 14809 14572 14924 14600
rect 14809 14569 14821 14572
rect 14763 14563 14821 14569
rect 14918 14560 14924 14572
rect 14976 14560 14982 14612
rect 17494 14600 17500 14612
rect 15732 14572 17500 14600
rect 12986 14492 12992 14544
rect 13044 14492 13050 14544
rect 13630 14492 13636 14544
rect 13688 14492 13694 14544
rect 14550 14492 14556 14544
rect 14608 14532 14614 14544
rect 15732 14532 15760 14572
rect 17494 14560 17500 14572
rect 17552 14560 17558 14612
rect 18046 14560 18052 14612
rect 18104 14600 18110 14612
rect 18233 14603 18291 14609
rect 18233 14600 18245 14603
rect 18104 14572 18245 14600
rect 18104 14560 18110 14572
rect 18233 14569 18245 14572
rect 18279 14569 18291 14603
rect 18233 14563 18291 14569
rect 18322 14560 18328 14612
rect 18380 14600 18386 14612
rect 18509 14603 18567 14609
rect 18509 14600 18521 14603
rect 18380 14572 18521 14600
rect 18380 14560 18386 14572
rect 18509 14569 18521 14572
rect 18555 14569 18567 14603
rect 18509 14563 18567 14569
rect 14608 14504 15760 14532
rect 16040 14504 17250 14532
rect 14608 14492 14614 14504
rect 12710 14424 12716 14476
rect 12768 14424 12774 14476
rect 16040 14464 16068 14504
rect 15212 14436 16068 14464
rect 18417 14467 18475 14473
rect 13722 14356 13728 14408
rect 13780 14396 13786 14408
rect 15212 14396 15240 14436
rect 18417 14433 18429 14467
rect 18463 14433 18475 14467
rect 18417 14427 18475 14433
rect 13780 14368 15240 14396
rect 13780 14356 13786 14368
rect 15286 14356 15292 14408
rect 15344 14396 15350 14408
rect 16482 14396 16488 14408
rect 15344 14368 16488 14396
rect 15344 14356 15350 14368
rect 16482 14356 16488 14368
rect 16540 14356 16546 14408
rect 16761 14399 16819 14405
rect 16761 14365 16773 14399
rect 16807 14396 16819 14399
rect 16850 14396 16856 14408
rect 16807 14368 16856 14396
rect 16807 14365 16819 14368
rect 16761 14359 16819 14365
rect 16850 14356 16856 14368
rect 16908 14356 16914 14408
rect 17126 14356 17132 14408
rect 17184 14396 17190 14408
rect 17770 14396 17776 14408
rect 17184 14368 17776 14396
rect 17184 14356 17190 14368
rect 17770 14356 17776 14368
rect 17828 14396 17834 14408
rect 18432 14396 18460 14427
rect 17828 14368 18460 14396
rect 17828 14356 17834 14368
rect 13998 14288 14004 14340
rect 14056 14328 14062 14340
rect 14056 14300 14780 14328
rect 14056 14288 14062 14300
rect 14752 14269 14780 14300
rect 31018 14288 31024 14340
rect 31076 14288 31082 14340
rect 14737 14263 14795 14269
rect 14737 14229 14749 14263
rect 14783 14229 14795 14263
rect 14737 14223 14795 14229
rect 14921 14263 14979 14269
rect 14921 14229 14933 14263
rect 14967 14260 14979 14263
rect 15010 14260 15016 14272
rect 14967 14232 15016 14260
rect 14967 14229 14979 14232
rect 14921 14223 14979 14229
rect 15010 14220 15016 14232
rect 15068 14220 15074 14272
rect 552 14170 31372 14192
rect 552 14118 3662 14170
rect 3714 14118 3726 14170
rect 3778 14118 3790 14170
rect 3842 14118 3854 14170
rect 3906 14118 3918 14170
rect 3970 14118 11436 14170
rect 11488 14118 11500 14170
rect 11552 14118 11564 14170
rect 11616 14118 11628 14170
rect 11680 14118 11692 14170
rect 11744 14118 19210 14170
rect 19262 14118 19274 14170
rect 19326 14118 19338 14170
rect 19390 14118 19402 14170
rect 19454 14118 19466 14170
rect 19518 14118 26984 14170
rect 27036 14118 27048 14170
rect 27100 14118 27112 14170
rect 27164 14118 27176 14170
rect 27228 14118 27240 14170
rect 27292 14118 31372 14170
rect 552 14096 31372 14118
rect 13541 14059 13599 14065
rect 13541 14025 13553 14059
rect 13587 14056 13599 14059
rect 13906 14056 13912 14068
rect 13587 14028 13912 14056
rect 13587 14025 13599 14028
rect 13541 14019 13599 14025
rect 13906 14016 13912 14028
rect 13964 14016 13970 14068
rect 16761 14059 16819 14065
rect 16761 14025 16773 14059
rect 16807 14056 16819 14059
rect 16850 14056 16856 14068
rect 16807 14028 16856 14056
rect 16807 14025 16819 14028
rect 16761 14019 16819 14025
rect 16850 14016 16856 14028
rect 16908 14016 16914 14068
rect 16942 14016 16948 14068
rect 17000 14016 17006 14068
rect 13814 13880 13820 13932
rect 13872 13880 13878 13932
rect 15010 13880 15016 13932
rect 15068 13880 15074 13932
rect 15286 13880 15292 13932
rect 15344 13880 15350 13932
rect 18046 13920 18052 13932
rect 17420 13892 18052 13920
rect 13832 13852 13860 13880
rect 17420 13861 17448 13892
rect 18046 13880 18052 13892
rect 18104 13880 18110 13932
rect 17221 13855 17279 13861
rect 17221 13852 17233 13855
rect 13832 13824 13938 13852
rect 16960 13824 17233 13852
rect 16960 13793 16988 13824
rect 17221 13821 17233 13824
rect 17267 13821 17279 13855
rect 17221 13815 17279 13821
rect 17405 13855 17463 13861
rect 17405 13821 17417 13855
rect 17451 13821 17463 13855
rect 17405 13815 17463 13821
rect 17589 13855 17647 13861
rect 17589 13821 17601 13855
rect 17635 13852 17647 13855
rect 17678 13852 17684 13864
rect 17635 13824 17684 13852
rect 17635 13821 17647 13824
rect 17589 13815 17647 13821
rect 17678 13812 17684 13824
rect 17736 13812 17742 13864
rect 16929 13787 16988 13793
rect 16929 13753 16941 13787
rect 16975 13756 16988 13787
rect 17129 13787 17187 13793
rect 16975 13753 16987 13756
rect 16929 13747 16987 13753
rect 17129 13753 17141 13787
rect 17175 13784 17187 13787
rect 17494 13784 17500 13796
rect 17175 13756 17500 13784
rect 17175 13753 17187 13756
rect 17129 13747 17187 13753
rect 17494 13744 17500 13756
rect 17552 13744 17558 13796
rect 552 13626 31372 13648
rect 552 13574 4322 13626
rect 4374 13574 4386 13626
rect 4438 13574 4450 13626
rect 4502 13574 4514 13626
rect 4566 13574 4578 13626
rect 4630 13574 12096 13626
rect 12148 13574 12160 13626
rect 12212 13574 12224 13626
rect 12276 13574 12288 13626
rect 12340 13574 12352 13626
rect 12404 13574 19870 13626
rect 19922 13574 19934 13626
rect 19986 13574 19998 13626
rect 20050 13574 20062 13626
rect 20114 13574 20126 13626
rect 20178 13574 27644 13626
rect 27696 13574 27708 13626
rect 27760 13574 27772 13626
rect 27824 13574 27836 13626
rect 27888 13574 27900 13626
rect 27952 13574 31372 13626
rect 552 13552 31372 13574
rect 552 13082 31372 13104
rect 552 13030 3662 13082
rect 3714 13030 3726 13082
rect 3778 13030 3790 13082
rect 3842 13030 3854 13082
rect 3906 13030 3918 13082
rect 3970 13030 11436 13082
rect 11488 13030 11500 13082
rect 11552 13030 11564 13082
rect 11616 13030 11628 13082
rect 11680 13030 11692 13082
rect 11744 13030 19210 13082
rect 19262 13030 19274 13082
rect 19326 13030 19338 13082
rect 19390 13030 19402 13082
rect 19454 13030 19466 13082
rect 19518 13030 26984 13082
rect 27036 13030 27048 13082
rect 27100 13030 27112 13082
rect 27164 13030 27176 13082
rect 27228 13030 27240 13082
rect 27292 13030 31372 13082
rect 552 13008 31372 13030
rect 552 12538 31372 12560
rect 552 12486 4322 12538
rect 4374 12486 4386 12538
rect 4438 12486 4450 12538
rect 4502 12486 4514 12538
rect 4566 12486 4578 12538
rect 4630 12486 12096 12538
rect 12148 12486 12160 12538
rect 12212 12486 12224 12538
rect 12276 12486 12288 12538
rect 12340 12486 12352 12538
rect 12404 12486 19870 12538
rect 19922 12486 19934 12538
rect 19986 12486 19998 12538
rect 20050 12486 20062 12538
rect 20114 12486 20126 12538
rect 20178 12486 27644 12538
rect 27696 12486 27708 12538
rect 27760 12486 27772 12538
rect 27824 12486 27836 12538
rect 27888 12486 27900 12538
rect 27952 12486 31372 12538
rect 552 12464 31372 12486
rect 552 11994 31372 12016
rect 552 11942 3662 11994
rect 3714 11942 3726 11994
rect 3778 11942 3790 11994
rect 3842 11942 3854 11994
rect 3906 11942 3918 11994
rect 3970 11942 11436 11994
rect 11488 11942 11500 11994
rect 11552 11942 11564 11994
rect 11616 11942 11628 11994
rect 11680 11942 11692 11994
rect 11744 11942 19210 11994
rect 19262 11942 19274 11994
rect 19326 11942 19338 11994
rect 19390 11942 19402 11994
rect 19454 11942 19466 11994
rect 19518 11942 26984 11994
rect 27036 11942 27048 11994
rect 27100 11942 27112 11994
rect 27164 11942 27176 11994
rect 27228 11942 27240 11994
rect 27292 11942 31372 11994
rect 552 11920 31372 11942
rect 552 11450 31372 11472
rect 552 11398 4322 11450
rect 4374 11398 4386 11450
rect 4438 11398 4450 11450
rect 4502 11398 4514 11450
rect 4566 11398 4578 11450
rect 4630 11398 12096 11450
rect 12148 11398 12160 11450
rect 12212 11398 12224 11450
rect 12276 11398 12288 11450
rect 12340 11398 12352 11450
rect 12404 11398 19870 11450
rect 19922 11398 19934 11450
rect 19986 11398 19998 11450
rect 20050 11398 20062 11450
rect 20114 11398 20126 11450
rect 20178 11398 27644 11450
rect 27696 11398 27708 11450
rect 27760 11398 27772 11450
rect 27824 11398 27836 11450
rect 27888 11398 27900 11450
rect 27952 11398 31372 11450
rect 552 11376 31372 11398
rect 552 10906 31372 10928
rect 552 10854 3662 10906
rect 3714 10854 3726 10906
rect 3778 10854 3790 10906
rect 3842 10854 3854 10906
rect 3906 10854 3918 10906
rect 3970 10854 11436 10906
rect 11488 10854 11500 10906
rect 11552 10854 11564 10906
rect 11616 10854 11628 10906
rect 11680 10854 11692 10906
rect 11744 10854 19210 10906
rect 19262 10854 19274 10906
rect 19326 10854 19338 10906
rect 19390 10854 19402 10906
rect 19454 10854 19466 10906
rect 19518 10854 26984 10906
rect 27036 10854 27048 10906
rect 27100 10854 27112 10906
rect 27164 10854 27176 10906
rect 27228 10854 27240 10906
rect 27292 10854 31372 10906
rect 552 10832 31372 10854
rect 552 10362 31372 10384
rect 552 10310 4322 10362
rect 4374 10310 4386 10362
rect 4438 10310 4450 10362
rect 4502 10310 4514 10362
rect 4566 10310 4578 10362
rect 4630 10310 12096 10362
rect 12148 10310 12160 10362
rect 12212 10310 12224 10362
rect 12276 10310 12288 10362
rect 12340 10310 12352 10362
rect 12404 10310 19870 10362
rect 19922 10310 19934 10362
rect 19986 10310 19998 10362
rect 20050 10310 20062 10362
rect 20114 10310 20126 10362
rect 20178 10310 27644 10362
rect 27696 10310 27708 10362
rect 27760 10310 27772 10362
rect 27824 10310 27836 10362
rect 27888 10310 27900 10362
rect 27952 10310 31372 10362
rect 552 10288 31372 10310
rect 552 9818 31372 9840
rect 552 9766 3662 9818
rect 3714 9766 3726 9818
rect 3778 9766 3790 9818
rect 3842 9766 3854 9818
rect 3906 9766 3918 9818
rect 3970 9766 11436 9818
rect 11488 9766 11500 9818
rect 11552 9766 11564 9818
rect 11616 9766 11628 9818
rect 11680 9766 11692 9818
rect 11744 9766 19210 9818
rect 19262 9766 19274 9818
rect 19326 9766 19338 9818
rect 19390 9766 19402 9818
rect 19454 9766 19466 9818
rect 19518 9766 26984 9818
rect 27036 9766 27048 9818
rect 27100 9766 27112 9818
rect 27164 9766 27176 9818
rect 27228 9766 27240 9818
rect 27292 9766 31372 9818
rect 552 9744 31372 9766
rect 552 9274 31372 9296
rect 552 9222 4322 9274
rect 4374 9222 4386 9274
rect 4438 9222 4450 9274
rect 4502 9222 4514 9274
rect 4566 9222 4578 9274
rect 4630 9222 12096 9274
rect 12148 9222 12160 9274
rect 12212 9222 12224 9274
rect 12276 9222 12288 9274
rect 12340 9222 12352 9274
rect 12404 9222 19870 9274
rect 19922 9222 19934 9274
rect 19986 9222 19998 9274
rect 20050 9222 20062 9274
rect 20114 9222 20126 9274
rect 20178 9222 27644 9274
rect 27696 9222 27708 9274
rect 27760 9222 27772 9274
rect 27824 9222 27836 9274
rect 27888 9222 27900 9274
rect 27952 9222 31372 9274
rect 552 9200 31372 9222
rect 552 8730 31372 8752
rect 552 8678 3662 8730
rect 3714 8678 3726 8730
rect 3778 8678 3790 8730
rect 3842 8678 3854 8730
rect 3906 8678 3918 8730
rect 3970 8678 11436 8730
rect 11488 8678 11500 8730
rect 11552 8678 11564 8730
rect 11616 8678 11628 8730
rect 11680 8678 11692 8730
rect 11744 8678 19210 8730
rect 19262 8678 19274 8730
rect 19326 8678 19338 8730
rect 19390 8678 19402 8730
rect 19454 8678 19466 8730
rect 19518 8678 26984 8730
rect 27036 8678 27048 8730
rect 27100 8678 27112 8730
rect 27164 8678 27176 8730
rect 27228 8678 27240 8730
rect 27292 8678 31372 8730
rect 552 8656 31372 8678
rect 552 8186 31372 8208
rect 552 8134 4322 8186
rect 4374 8134 4386 8186
rect 4438 8134 4450 8186
rect 4502 8134 4514 8186
rect 4566 8134 4578 8186
rect 4630 8134 12096 8186
rect 12148 8134 12160 8186
rect 12212 8134 12224 8186
rect 12276 8134 12288 8186
rect 12340 8134 12352 8186
rect 12404 8134 19870 8186
rect 19922 8134 19934 8186
rect 19986 8134 19998 8186
rect 20050 8134 20062 8186
rect 20114 8134 20126 8186
rect 20178 8134 27644 8186
rect 27696 8134 27708 8186
rect 27760 8134 27772 8186
rect 27824 8134 27836 8186
rect 27888 8134 27900 8186
rect 27952 8134 31372 8186
rect 552 8112 31372 8134
rect 552 7642 31372 7664
rect 552 7590 3662 7642
rect 3714 7590 3726 7642
rect 3778 7590 3790 7642
rect 3842 7590 3854 7642
rect 3906 7590 3918 7642
rect 3970 7590 11436 7642
rect 11488 7590 11500 7642
rect 11552 7590 11564 7642
rect 11616 7590 11628 7642
rect 11680 7590 11692 7642
rect 11744 7590 19210 7642
rect 19262 7590 19274 7642
rect 19326 7590 19338 7642
rect 19390 7590 19402 7642
rect 19454 7590 19466 7642
rect 19518 7590 26984 7642
rect 27036 7590 27048 7642
rect 27100 7590 27112 7642
rect 27164 7590 27176 7642
rect 27228 7590 27240 7642
rect 27292 7590 31372 7642
rect 552 7568 31372 7590
rect 552 7098 31372 7120
rect 552 7046 4322 7098
rect 4374 7046 4386 7098
rect 4438 7046 4450 7098
rect 4502 7046 4514 7098
rect 4566 7046 4578 7098
rect 4630 7046 12096 7098
rect 12148 7046 12160 7098
rect 12212 7046 12224 7098
rect 12276 7046 12288 7098
rect 12340 7046 12352 7098
rect 12404 7046 19870 7098
rect 19922 7046 19934 7098
rect 19986 7046 19998 7098
rect 20050 7046 20062 7098
rect 20114 7046 20126 7098
rect 20178 7046 27644 7098
rect 27696 7046 27708 7098
rect 27760 7046 27772 7098
rect 27824 7046 27836 7098
rect 27888 7046 27900 7098
rect 27952 7046 31372 7098
rect 552 7024 31372 7046
rect 552 6554 31372 6576
rect 552 6502 3662 6554
rect 3714 6502 3726 6554
rect 3778 6502 3790 6554
rect 3842 6502 3854 6554
rect 3906 6502 3918 6554
rect 3970 6502 11436 6554
rect 11488 6502 11500 6554
rect 11552 6502 11564 6554
rect 11616 6502 11628 6554
rect 11680 6502 11692 6554
rect 11744 6502 19210 6554
rect 19262 6502 19274 6554
rect 19326 6502 19338 6554
rect 19390 6502 19402 6554
rect 19454 6502 19466 6554
rect 19518 6502 26984 6554
rect 27036 6502 27048 6554
rect 27100 6502 27112 6554
rect 27164 6502 27176 6554
rect 27228 6502 27240 6554
rect 27292 6502 31372 6554
rect 552 6480 31372 6502
rect 552 6010 31372 6032
rect 552 5958 4322 6010
rect 4374 5958 4386 6010
rect 4438 5958 4450 6010
rect 4502 5958 4514 6010
rect 4566 5958 4578 6010
rect 4630 5958 12096 6010
rect 12148 5958 12160 6010
rect 12212 5958 12224 6010
rect 12276 5958 12288 6010
rect 12340 5958 12352 6010
rect 12404 5958 19870 6010
rect 19922 5958 19934 6010
rect 19986 5958 19998 6010
rect 20050 5958 20062 6010
rect 20114 5958 20126 6010
rect 20178 5958 27644 6010
rect 27696 5958 27708 6010
rect 27760 5958 27772 6010
rect 27824 5958 27836 6010
rect 27888 5958 27900 6010
rect 27952 5958 31372 6010
rect 552 5936 31372 5958
rect 552 5466 31372 5488
rect 552 5414 3662 5466
rect 3714 5414 3726 5466
rect 3778 5414 3790 5466
rect 3842 5414 3854 5466
rect 3906 5414 3918 5466
rect 3970 5414 11436 5466
rect 11488 5414 11500 5466
rect 11552 5414 11564 5466
rect 11616 5414 11628 5466
rect 11680 5414 11692 5466
rect 11744 5414 19210 5466
rect 19262 5414 19274 5466
rect 19326 5414 19338 5466
rect 19390 5414 19402 5466
rect 19454 5414 19466 5466
rect 19518 5414 26984 5466
rect 27036 5414 27048 5466
rect 27100 5414 27112 5466
rect 27164 5414 27176 5466
rect 27228 5414 27240 5466
rect 27292 5414 31372 5466
rect 552 5392 31372 5414
rect 552 4922 31372 4944
rect 552 4870 4322 4922
rect 4374 4870 4386 4922
rect 4438 4870 4450 4922
rect 4502 4870 4514 4922
rect 4566 4870 4578 4922
rect 4630 4870 12096 4922
rect 12148 4870 12160 4922
rect 12212 4870 12224 4922
rect 12276 4870 12288 4922
rect 12340 4870 12352 4922
rect 12404 4870 19870 4922
rect 19922 4870 19934 4922
rect 19986 4870 19998 4922
rect 20050 4870 20062 4922
rect 20114 4870 20126 4922
rect 20178 4870 27644 4922
rect 27696 4870 27708 4922
rect 27760 4870 27772 4922
rect 27824 4870 27836 4922
rect 27888 4870 27900 4922
rect 27952 4870 31372 4922
rect 552 4848 31372 4870
rect 552 4378 31372 4400
rect 552 4326 3662 4378
rect 3714 4326 3726 4378
rect 3778 4326 3790 4378
rect 3842 4326 3854 4378
rect 3906 4326 3918 4378
rect 3970 4326 11436 4378
rect 11488 4326 11500 4378
rect 11552 4326 11564 4378
rect 11616 4326 11628 4378
rect 11680 4326 11692 4378
rect 11744 4326 19210 4378
rect 19262 4326 19274 4378
rect 19326 4326 19338 4378
rect 19390 4326 19402 4378
rect 19454 4326 19466 4378
rect 19518 4326 26984 4378
rect 27036 4326 27048 4378
rect 27100 4326 27112 4378
rect 27164 4326 27176 4378
rect 27228 4326 27240 4378
rect 27292 4326 31372 4378
rect 552 4304 31372 4326
rect 552 3834 31372 3856
rect 552 3782 4322 3834
rect 4374 3782 4386 3834
rect 4438 3782 4450 3834
rect 4502 3782 4514 3834
rect 4566 3782 4578 3834
rect 4630 3782 12096 3834
rect 12148 3782 12160 3834
rect 12212 3782 12224 3834
rect 12276 3782 12288 3834
rect 12340 3782 12352 3834
rect 12404 3782 19870 3834
rect 19922 3782 19934 3834
rect 19986 3782 19998 3834
rect 20050 3782 20062 3834
rect 20114 3782 20126 3834
rect 20178 3782 27644 3834
rect 27696 3782 27708 3834
rect 27760 3782 27772 3834
rect 27824 3782 27836 3834
rect 27888 3782 27900 3834
rect 27952 3782 31372 3834
rect 552 3760 31372 3782
rect 552 3290 31372 3312
rect 552 3238 3662 3290
rect 3714 3238 3726 3290
rect 3778 3238 3790 3290
rect 3842 3238 3854 3290
rect 3906 3238 3918 3290
rect 3970 3238 11436 3290
rect 11488 3238 11500 3290
rect 11552 3238 11564 3290
rect 11616 3238 11628 3290
rect 11680 3238 11692 3290
rect 11744 3238 19210 3290
rect 19262 3238 19274 3290
rect 19326 3238 19338 3290
rect 19390 3238 19402 3290
rect 19454 3238 19466 3290
rect 19518 3238 26984 3290
rect 27036 3238 27048 3290
rect 27100 3238 27112 3290
rect 27164 3238 27176 3290
rect 27228 3238 27240 3290
rect 27292 3238 31372 3290
rect 552 3216 31372 3238
rect 552 2746 31372 2768
rect 552 2694 4322 2746
rect 4374 2694 4386 2746
rect 4438 2694 4450 2746
rect 4502 2694 4514 2746
rect 4566 2694 4578 2746
rect 4630 2694 12096 2746
rect 12148 2694 12160 2746
rect 12212 2694 12224 2746
rect 12276 2694 12288 2746
rect 12340 2694 12352 2746
rect 12404 2694 19870 2746
rect 19922 2694 19934 2746
rect 19986 2694 19998 2746
rect 20050 2694 20062 2746
rect 20114 2694 20126 2746
rect 20178 2694 27644 2746
rect 27696 2694 27708 2746
rect 27760 2694 27772 2746
rect 27824 2694 27836 2746
rect 27888 2694 27900 2746
rect 27952 2694 31372 2746
rect 552 2672 31372 2694
rect 552 2202 31372 2224
rect 552 2150 3662 2202
rect 3714 2150 3726 2202
rect 3778 2150 3790 2202
rect 3842 2150 3854 2202
rect 3906 2150 3918 2202
rect 3970 2150 11436 2202
rect 11488 2150 11500 2202
rect 11552 2150 11564 2202
rect 11616 2150 11628 2202
rect 11680 2150 11692 2202
rect 11744 2150 19210 2202
rect 19262 2150 19274 2202
rect 19326 2150 19338 2202
rect 19390 2150 19402 2202
rect 19454 2150 19466 2202
rect 19518 2150 26984 2202
rect 27036 2150 27048 2202
rect 27100 2150 27112 2202
rect 27164 2150 27176 2202
rect 27228 2150 27240 2202
rect 27292 2150 31372 2202
rect 552 2128 31372 2150
rect 552 1658 31372 1680
rect 552 1606 4322 1658
rect 4374 1606 4386 1658
rect 4438 1606 4450 1658
rect 4502 1606 4514 1658
rect 4566 1606 4578 1658
rect 4630 1606 12096 1658
rect 12148 1606 12160 1658
rect 12212 1606 12224 1658
rect 12276 1606 12288 1658
rect 12340 1606 12352 1658
rect 12404 1606 19870 1658
rect 19922 1606 19934 1658
rect 19986 1606 19998 1658
rect 20050 1606 20062 1658
rect 20114 1606 20126 1658
rect 20178 1606 27644 1658
rect 27696 1606 27708 1658
rect 27760 1606 27772 1658
rect 27824 1606 27836 1658
rect 27888 1606 27900 1658
rect 27952 1606 31372 1658
rect 552 1584 31372 1606
rect 552 1114 31372 1136
rect 552 1062 3662 1114
rect 3714 1062 3726 1114
rect 3778 1062 3790 1114
rect 3842 1062 3854 1114
rect 3906 1062 3918 1114
rect 3970 1062 11436 1114
rect 11488 1062 11500 1114
rect 11552 1062 11564 1114
rect 11616 1062 11628 1114
rect 11680 1062 11692 1114
rect 11744 1062 19210 1114
rect 19262 1062 19274 1114
rect 19326 1062 19338 1114
rect 19390 1062 19402 1114
rect 19454 1062 19466 1114
rect 19518 1062 26984 1114
rect 27036 1062 27048 1114
rect 27100 1062 27112 1114
rect 27164 1062 27176 1114
rect 27228 1062 27240 1114
rect 27292 1062 31372 1114
rect 552 1040 31372 1062
rect 17034 960 17040 1012
rect 17092 960 17098 1012
rect 16114 892 16120 944
rect 16172 932 16178 944
rect 16758 932 16764 944
rect 16172 904 16764 932
rect 16172 892 16178 904
rect 16758 892 16764 904
rect 16816 892 16822 944
rect 7098 756 7104 808
rect 7156 796 7162 808
rect 7193 799 7251 805
rect 7193 796 7205 799
rect 7156 768 7205 796
rect 7156 756 7162 768
rect 7193 765 7205 768
rect 7239 765 7251 799
rect 7193 759 7251 765
rect 9030 756 9036 808
rect 9088 796 9094 808
rect 9125 799 9183 805
rect 9125 796 9137 799
rect 9088 768 9137 796
rect 9088 756 9094 768
rect 9125 765 9137 768
rect 9171 765 9183 799
rect 9125 759 9183 765
rect 11606 756 11612 808
rect 11664 796 11670 808
rect 11701 799 11759 805
rect 11701 796 11713 799
rect 11664 768 11713 796
rect 11664 756 11670 768
rect 11701 765 11713 768
rect 11747 765 11759 799
rect 11701 759 11759 765
rect 12345 799 12403 805
rect 12345 765 12357 799
rect 12391 796 12403 799
rect 12434 796 12440 808
rect 12391 768 12440 796
rect 12391 765 12403 768
rect 12345 759 12403 765
rect 12434 756 12440 768
rect 12492 756 12498 808
rect 12894 756 12900 808
rect 12952 796 12958 808
rect 12989 799 13047 805
rect 12989 796 13001 799
rect 12952 768 13001 796
rect 12952 756 12958 768
rect 12989 765 13001 768
rect 13035 765 13047 799
rect 12989 759 13047 765
rect 13538 756 13544 808
rect 13596 796 13602 808
rect 13633 799 13691 805
rect 13633 796 13645 799
rect 13596 768 13645 796
rect 13596 756 13602 768
rect 13633 765 13645 768
rect 13679 765 13691 799
rect 13633 759 13691 765
rect 14182 756 14188 808
rect 14240 796 14246 808
rect 14277 799 14335 805
rect 14277 796 14289 799
rect 14240 768 14289 796
rect 14240 756 14246 768
rect 14277 765 14289 768
rect 14323 765 14335 799
rect 14277 759 14335 765
rect 14826 756 14832 808
rect 14884 796 14890 808
rect 14921 799 14979 805
rect 14921 796 14933 799
rect 14884 768 14933 796
rect 14884 756 14890 768
rect 14921 765 14933 768
rect 14967 765 14979 799
rect 14921 759 14979 765
rect 15470 756 15476 808
rect 15528 796 15534 808
rect 15565 799 15623 805
rect 15565 796 15577 799
rect 15528 768 15577 796
rect 15528 756 15534 768
rect 15565 765 15577 768
rect 15611 765 15623 799
rect 15565 759 15623 765
rect 16758 756 16764 808
rect 16816 796 16822 808
rect 16853 799 16911 805
rect 16853 796 16865 799
rect 16816 768 16865 796
rect 16816 756 16822 768
rect 16853 765 16865 768
rect 16899 765 16911 799
rect 16853 759 16911 765
rect 17402 756 17408 808
rect 17460 796 17466 808
rect 17497 799 17555 805
rect 17497 796 17509 799
rect 17460 768 17509 796
rect 17460 756 17466 768
rect 17497 765 17509 768
rect 17543 765 17555 799
rect 17497 759 17555 765
rect 18046 756 18052 808
rect 18104 796 18110 808
rect 18141 799 18199 805
rect 18141 796 18153 799
rect 18104 768 18153 796
rect 18104 756 18110 768
rect 18141 765 18153 768
rect 18187 765 18199 799
rect 18141 759 18199 765
rect 18690 756 18696 808
rect 18748 796 18754 808
rect 18785 799 18843 805
rect 18785 796 18797 799
rect 18748 768 18797 796
rect 18748 756 18754 768
rect 18785 765 18797 768
rect 18831 765 18843 799
rect 18785 759 18843 765
rect 19794 756 19800 808
rect 19852 796 19858 808
rect 20073 799 20131 805
rect 20073 796 20085 799
rect 19852 768 20085 796
rect 19852 756 19858 768
rect 20073 765 20085 768
rect 20119 765 20131 799
rect 20073 759 20131 765
rect 552 570 31372 592
rect 552 518 4322 570
rect 4374 518 4386 570
rect 4438 518 4450 570
rect 4502 518 4514 570
rect 4566 518 4578 570
rect 4630 518 12096 570
rect 12148 518 12160 570
rect 12212 518 12224 570
rect 12276 518 12288 570
rect 12340 518 12352 570
rect 12404 518 19870 570
rect 19922 518 19934 570
rect 19986 518 19998 570
rect 20050 518 20062 570
rect 20114 518 20126 570
rect 20178 518 27644 570
rect 27696 518 27708 570
rect 27760 518 27772 570
rect 27824 518 27836 570
rect 27888 518 27900 570
rect 27952 518 31372 570
rect 552 496 31372 518
rect 12158 416 12164 468
rect 12216 456 12222 468
rect 12434 456 12440 468
rect 12216 428 12440 456
rect 12216 416 12222 428
rect 12434 416 12440 428
rect 12492 416 12498 468
<< via1 >>
rect 4322 19014 4374 19066
rect 4386 19014 4438 19066
rect 4450 19014 4502 19066
rect 4514 19014 4566 19066
rect 4578 19014 4630 19066
rect 12096 19014 12148 19066
rect 12160 19014 12212 19066
rect 12224 19014 12276 19066
rect 12288 19014 12340 19066
rect 12352 19014 12404 19066
rect 19870 19014 19922 19066
rect 19934 19014 19986 19066
rect 19998 19014 20050 19066
rect 20062 19014 20114 19066
rect 20126 19014 20178 19066
rect 27644 19014 27696 19066
rect 27708 19014 27760 19066
rect 27772 19014 27824 19066
rect 27836 19014 27888 19066
rect 27900 19014 27952 19066
rect 14832 18912 14884 18964
rect 16120 18912 16172 18964
rect 10324 18776 10376 18828
rect 11980 18776 12032 18828
rect 12900 18776 12952 18828
rect 13544 18776 13596 18828
rect 14188 18776 14240 18828
rect 17316 18776 17368 18828
rect 15292 18708 15344 18760
rect 22560 18776 22612 18828
rect 16764 18640 16816 18692
rect 848 18615 900 18624
rect 848 18581 857 18615
rect 857 18581 891 18615
rect 891 18581 900 18615
rect 848 18572 900 18581
rect 14372 18572 14424 18624
rect 15200 18615 15252 18624
rect 15200 18581 15209 18615
rect 15209 18581 15243 18615
rect 15243 18581 15252 18615
rect 15200 18572 15252 18581
rect 15384 18572 15436 18624
rect 18236 18615 18288 18624
rect 18236 18581 18245 18615
rect 18245 18581 18279 18615
rect 18279 18581 18288 18615
rect 18236 18572 18288 18581
rect 3662 18470 3714 18522
rect 3726 18470 3778 18522
rect 3790 18470 3842 18522
rect 3854 18470 3906 18522
rect 3918 18470 3970 18522
rect 11436 18470 11488 18522
rect 11500 18470 11552 18522
rect 11564 18470 11616 18522
rect 11628 18470 11680 18522
rect 11692 18470 11744 18522
rect 19210 18470 19262 18522
rect 19274 18470 19326 18522
rect 19338 18470 19390 18522
rect 19402 18470 19454 18522
rect 19466 18470 19518 18522
rect 26984 18470 27036 18522
rect 27048 18470 27100 18522
rect 27112 18470 27164 18522
rect 27176 18470 27228 18522
rect 27240 18470 27292 18522
rect 15292 18411 15344 18420
rect 15292 18377 15301 18411
rect 15301 18377 15335 18411
rect 15335 18377 15344 18411
rect 15292 18368 15344 18377
rect 17316 18368 17368 18420
rect 17500 18368 17552 18420
rect 14188 18232 14240 18284
rect 16396 18232 16448 18284
rect 17132 18232 17184 18284
rect 12716 18164 12768 18216
rect 15844 18207 15896 18216
rect 15844 18173 15853 18207
rect 15853 18173 15887 18207
rect 15887 18173 15896 18207
rect 15844 18164 15896 18173
rect 16764 18164 16816 18216
rect 13636 18028 13688 18080
rect 17684 18028 17736 18080
rect 17776 18071 17828 18080
rect 17776 18037 17785 18071
rect 17785 18037 17819 18071
rect 17819 18037 17828 18071
rect 17776 18028 17828 18037
rect 4322 17926 4374 17978
rect 4386 17926 4438 17978
rect 4450 17926 4502 17978
rect 4514 17926 4566 17978
rect 4578 17926 4630 17978
rect 12096 17926 12148 17978
rect 12160 17926 12212 17978
rect 12224 17926 12276 17978
rect 12288 17926 12340 17978
rect 12352 17926 12404 17978
rect 19870 17926 19922 17978
rect 19934 17926 19986 17978
rect 19998 17926 20050 17978
rect 20062 17926 20114 17978
rect 20126 17926 20178 17978
rect 27644 17926 27696 17978
rect 27708 17926 27760 17978
rect 27772 17926 27824 17978
rect 27836 17926 27888 17978
rect 27900 17926 27952 17978
rect 13636 17688 13688 17740
rect 14740 17756 14792 17808
rect 15200 17756 15252 17808
rect 15844 17824 15896 17876
rect 18236 17824 18288 17876
rect 14648 17731 14700 17740
rect 14648 17697 14657 17731
rect 14657 17697 14691 17731
rect 14691 17697 14700 17731
rect 14648 17688 14700 17697
rect 12532 17663 12584 17672
rect 12532 17629 12541 17663
rect 12541 17629 12575 17663
rect 12575 17629 12584 17663
rect 12532 17620 12584 17629
rect 14372 17663 14424 17672
rect 14372 17629 14381 17663
rect 14381 17629 14415 17663
rect 14415 17629 14424 17663
rect 14372 17620 14424 17629
rect 14648 17552 14700 17604
rect 12716 17484 12768 17536
rect 14004 17527 14056 17536
rect 14004 17493 14013 17527
rect 14013 17493 14047 17527
rect 14047 17493 14056 17527
rect 14004 17484 14056 17493
rect 14188 17484 14240 17536
rect 15016 17731 15068 17740
rect 15016 17697 15025 17731
rect 15025 17697 15059 17731
rect 15059 17697 15068 17731
rect 15016 17688 15068 17697
rect 16856 17688 16908 17740
rect 15292 17663 15344 17672
rect 15292 17629 15301 17663
rect 15301 17629 15335 17663
rect 15335 17629 15344 17663
rect 15292 17620 15344 17629
rect 16304 17620 16356 17672
rect 17960 17756 18012 17808
rect 19064 17756 19116 17808
rect 17132 17688 17184 17740
rect 17316 17620 17368 17672
rect 17592 17620 17644 17672
rect 16764 17484 16816 17536
rect 17408 17527 17460 17536
rect 17408 17493 17417 17527
rect 17417 17493 17451 17527
rect 17451 17493 17460 17527
rect 17408 17484 17460 17493
rect 3662 17382 3714 17434
rect 3726 17382 3778 17434
rect 3790 17382 3842 17434
rect 3854 17382 3906 17434
rect 3918 17382 3970 17434
rect 11436 17382 11488 17434
rect 11500 17382 11552 17434
rect 11564 17382 11616 17434
rect 11628 17382 11680 17434
rect 11692 17382 11744 17434
rect 19210 17382 19262 17434
rect 19274 17382 19326 17434
rect 19338 17382 19390 17434
rect 19402 17382 19454 17434
rect 19466 17382 19518 17434
rect 26984 17382 27036 17434
rect 27048 17382 27100 17434
rect 27112 17382 27164 17434
rect 27176 17382 27228 17434
rect 27240 17382 27292 17434
rect 14648 17280 14700 17332
rect 15108 17280 15160 17332
rect 16304 17280 16356 17332
rect 16764 17323 16816 17332
rect 16764 17289 16773 17323
rect 16773 17289 16807 17323
rect 16807 17289 16816 17323
rect 16764 17280 16816 17289
rect 16856 17323 16908 17332
rect 16856 17289 16865 17323
rect 16865 17289 16899 17323
rect 16899 17289 16908 17323
rect 16856 17280 16908 17289
rect 17592 17323 17644 17332
rect 17592 17289 17601 17323
rect 17601 17289 17635 17323
rect 17635 17289 17644 17323
rect 17592 17280 17644 17289
rect 17776 17323 17828 17332
rect 17776 17289 17785 17323
rect 17785 17289 17819 17323
rect 17819 17289 17828 17323
rect 17776 17280 17828 17289
rect 12716 17212 12768 17264
rect 13636 17144 13688 17196
rect 13728 17119 13780 17128
rect 13728 17085 13737 17119
rect 13737 17085 13771 17119
rect 13771 17085 13780 17119
rect 13728 17076 13780 17085
rect 14004 17119 14056 17128
rect 14004 17085 14013 17119
rect 14013 17085 14047 17119
rect 14047 17085 14056 17119
rect 14004 17076 14056 17085
rect 12716 17008 12768 17060
rect 15292 17187 15344 17196
rect 15292 17153 15301 17187
rect 15301 17153 15335 17187
rect 15335 17153 15344 17187
rect 15292 17144 15344 17153
rect 18328 17144 18380 17196
rect 17960 17076 18012 17128
rect 13820 16983 13872 16992
rect 13820 16949 13829 16983
rect 13829 16949 13863 16983
rect 13863 16949 13872 16983
rect 13820 16940 13872 16949
rect 14188 16983 14240 16992
rect 14188 16949 14197 16983
rect 14197 16949 14231 16983
rect 14231 16949 14240 16983
rect 14188 16940 14240 16949
rect 14832 16983 14884 16992
rect 14832 16949 14841 16983
rect 14841 16949 14875 16983
rect 14875 16949 14884 16983
rect 14832 16940 14884 16949
rect 15384 17008 15436 17060
rect 17316 17008 17368 17060
rect 17408 17008 17460 17060
rect 17684 17008 17736 17060
rect 16672 16940 16724 16992
rect 17500 16940 17552 16992
rect 4322 16838 4374 16890
rect 4386 16838 4438 16890
rect 4450 16838 4502 16890
rect 4514 16838 4566 16890
rect 4578 16838 4630 16890
rect 12096 16838 12148 16890
rect 12160 16838 12212 16890
rect 12224 16838 12276 16890
rect 12288 16838 12340 16890
rect 12352 16838 12404 16890
rect 19870 16838 19922 16890
rect 19934 16838 19986 16890
rect 19998 16838 20050 16890
rect 20062 16838 20114 16890
rect 20126 16838 20178 16890
rect 27644 16838 27696 16890
rect 27708 16838 27760 16890
rect 27772 16838 27824 16890
rect 27836 16838 27888 16890
rect 27900 16838 27952 16890
rect 14188 16736 14240 16788
rect 15476 16736 15528 16788
rect 16672 16668 16724 16720
rect 12532 16600 12584 16652
rect 14832 16643 14884 16652
rect 14832 16609 14841 16643
rect 14841 16609 14875 16643
rect 14875 16609 14884 16643
rect 14832 16600 14884 16609
rect 15200 16600 15252 16652
rect 15568 16643 15620 16652
rect 15568 16609 15577 16643
rect 15577 16609 15611 16643
rect 15611 16609 15620 16643
rect 15568 16600 15620 16609
rect 12716 16575 12768 16584
rect 12716 16541 12725 16575
rect 12725 16541 12759 16575
rect 12759 16541 12768 16575
rect 12716 16532 12768 16541
rect 16580 16600 16632 16652
rect 17132 16668 17184 16720
rect 17316 16668 17368 16720
rect 17040 16643 17092 16652
rect 17040 16609 17049 16643
rect 17049 16609 17083 16643
rect 17083 16609 17092 16643
rect 17040 16600 17092 16609
rect 17224 16643 17276 16652
rect 17224 16609 17233 16643
rect 17233 16609 17267 16643
rect 17267 16609 17276 16643
rect 17224 16600 17276 16609
rect 19156 16643 19208 16652
rect 19156 16609 19165 16643
rect 19165 16609 19199 16643
rect 19199 16609 19208 16643
rect 19156 16600 19208 16609
rect 18880 16575 18932 16584
rect 18880 16541 18889 16575
rect 18889 16541 18923 16575
rect 18923 16541 18932 16575
rect 18880 16532 18932 16541
rect 14004 16464 14056 16516
rect 15568 16464 15620 16516
rect 16948 16464 17000 16516
rect 19156 16464 19208 16516
rect 15844 16396 15896 16448
rect 16672 16439 16724 16448
rect 16672 16405 16681 16439
rect 16681 16405 16715 16439
rect 16715 16405 16724 16439
rect 16672 16396 16724 16405
rect 17040 16396 17092 16448
rect 3662 16294 3714 16346
rect 3726 16294 3778 16346
rect 3790 16294 3842 16346
rect 3854 16294 3906 16346
rect 3918 16294 3970 16346
rect 11436 16294 11488 16346
rect 11500 16294 11552 16346
rect 11564 16294 11616 16346
rect 11628 16294 11680 16346
rect 11692 16294 11744 16346
rect 19210 16294 19262 16346
rect 19274 16294 19326 16346
rect 19338 16294 19390 16346
rect 19402 16294 19454 16346
rect 19466 16294 19518 16346
rect 26984 16294 27036 16346
rect 27048 16294 27100 16346
rect 27112 16294 27164 16346
rect 27176 16294 27228 16346
rect 27240 16294 27292 16346
rect 12808 16192 12860 16244
rect 14556 16192 14608 16244
rect 15476 16235 15528 16244
rect 15476 16201 15485 16235
rect 15485 16201 15519 16235
rect 15519 16201 15528 16235
rect 15476 16192 15528 16201
rect 14004 16124 14056 16176
rect 14372 16056 14424 16108
rect 15752 16056 15804 16108
rect 18236 16124 18288 16176
rect 19340 16192 19392 16244
rect 12992 15988 13044 16040
rect 13728 16031 13780 16040
rect 13728 15997 13737 16031
rect 13737 15997 13771 16031
rect 13771 15997 13780 16031
rect 13728 15988 13780 15997
rect 13820 16031 13872 16040
rect 13820 15997 13829 16031
rect 13829 15997 13863 16031
rect 13863 15997 13872 16031
rect 13820 15988 13872 15997
rect 14004 16031 14056 16040
rect 14004 15997 14013 16031
rect 14013 15997 14047 16031
rect 14047 15997 14056 16031
rect 14004 15988 14056 15997
rect 17040 15988 17092 16040
rect 17224 15988 17276 16040
rect 14372 15920 14424 15972
rect 16764 15963 16816 15972
rect 16764 15929 16773 15963
rect 16773 15929 16807 15963
rect 16807 15929 16816 15963
rect 16764 15920 16816 15929
rect 18052 15920 18104 15972
rect 18328 15963 18380 15972
rect 12532 15852 12584 15904
rect 16856 15852 16908 15904
rect 17132 15852 17184 15904
rect 17316 15895 17368 15904
rect 17316 15861 17325 15895
rect 17325 15861 17359 15895
rect 17359 15861 17368 15895
rect 17316 15852 17368 15861
rect 17408 15895 17460 15904
rect 17408 15861 17417 15895
rect 17417 15861 17451 15895
rect 17451 15861 17460 15895
rect 17408 15852 17460 15861
rect 17592 15852 17644 15904
rect 18328 15929 18355 15963
rect 18355 15929 18380 15963
rect 18328 15920 18380 15929
rect 4322 15750 4374 15802
rect 4386 15750 4438 15802
rect 4450 15750 4502 15802
rect 4514 15750 4566 15802
rect 4578 15750 4630 15802
rect 12096 15750 12148 15802
rect 12160 15750 12212 15802
rect 12224 15750 12276 15802
rect 12288 15750 12340 15802
rect 12352 15750 12404 15802
rect 19870 15750 19922 15802
rect 19934 15750 19986 15802
rect 19998 15750 20050 15802
rect 20062 15750 20114 15802
rect 20126 15750 20178 15802
rect 27644 15750 27696 15802
rect 27708 15750 27760 15802
rect 27772 15750 27824 15802
rect 27836 15750 27888 15802
rect 27900 15750 27952 15802
rect 14004 15691 14056 15700
rect 14004 15657 14013 15691
rect 14013 15657 14047 15691
rect 14047 15657 14056 15691
rect 14004 15648 14056 15657
rect 14096 15648 14148 15700
rect 14740 15648 14792 15700
rect 12532 15623 12584 15632
rect 12532 15589 12541 15623
rect 12541 15589 12575 15623
rect 12575 15589 12584 15623
rect 12532 15580 12584 15589
rect 13636 15512 13688 15564
rect 13820 15512 13872 15564
rect 12992 15444 13044 15496
rect 14372 15555 14424 15564
rect 14372 15521 14381 15555
rect 14381 15521 14415 15555
rect 14415 15521 14424 15555
rect 14372 15512 14424 15521
rect 14464 15512 14516 15564
rect 14924 15555 14976 15564
rect 14924 15521 14933 15555
rect 14933 15521 14967 15555
rect 14967 15521 14976 15555
rect 14924 15512 14976 15521
rect 15844 15623 15896 15632
rect 15844 15589 15853 15623
rect 15853 15589 15887 15623
rect 15887 15589 15896 15623
rect 15844 15580 15896 15589
rect 15476 15512 15528 15564
rect 15752 15555 15804 15564
rect 15752 15521 15761 15555
rect 15761 15521 15795 15555
rect 15795 15521 15804 15555
rect 15752 15512 15804 15521
rect 15568 15444 15620 15496
rect 15936 15555 15988 15564
rect 15936 15521 15945 15555
rect 15945 15521 15979 15555
rect 15979 15521 15988 15555
rect 15936 15512 15988 15521
rect 16488 15555 16540 15564
rect 16488 15521 16497 15555
rect 16497 15521 16531 15555
rect 16531 15521 16540 15555
rect 16488 15512 16540 15521
rect 16948 15648 17000 15700
rect 17500 15648 17552 15700
rect 18880 15648 18932 15700
rect 19340 15691 19392 15700
rect 19340 15657 19349 15691
rect 19349 15657 19383 15691
rect 19383 15657 19392 15691
rect 19340 15648 19392 15657
rect 16672 15512 16724 15564
rect 17132 15555 17184 15564
rect 17132 15521 17141 15555
rect 17141 15521 17175 15555
rect 17175 15521 17184 15555
rect 17132 15512 17184 15521
rect 17408 15512 17460 15564
rect 17960 15580 18012 15632
rect 18328 15580 18380 15632
rect 13912 15376 13964 15428
rect 14924 15376 14976 15428
rect 15200 15376 15252 15428
rect 16488 15376 16540 15428
rect 12716 15308 12768 15360
rect 14740 15351 14792 15360
rect 14740 15317 14749 15351
rect 14749 15317 14783 15351
rect 14783 15317 14792 15351
rect 14740 15308 14792 15317
rect 17040 15308 17092 15360
rect 17868 15487 17920 15496
rect 17868 15453 17877 15487
rect 17877 15453 17911 15487
rect 17911 15453 17920 15487
rect 17868 15444 17920 15453
rect 19064 15308 19116 15360
rect 3662 15206 3714 15258
rect 3726 15206 3778 15258
rect 3790 15206 3842 15258
rect 3854 15206 3906 15258
rect 3918 15206 3970 15258
rect 11436 15206 11488 15258
rect 11500 15206 11552 15258
rect 11564 15206 11616 15258
rect 11628 15206 11680 15258
rect 11692 15206 11744 15258
rect 19210 15206 19262 15258
rect 19274 15206 19326 15258
rect 19338 15206 19390 15258
rect 19402 15206 19454 15258
rect 19466 15206 19518 15258
rect 26984 15206 27036 15258
rect 27048 15206 27100 15258
rect 27112 15206 27164 15258
rect 27176 15206 27228 15258
rect 27240 15206 27292 15258
rect 12624 15104 12676 15156
rect 14740 15104 14792 15156
rect 15936 15104 15988 15156
rect 17040 15104 17092 15156
rect 17500 15147 17552 15156
rect 17500 15113 17509 15147
rect 17509 15113 17543 15147
rect 17543 15113 17552 15147
rect 17500 15104 17552 15113
rect 17868 15104 17920 15156
rect 12532 15036 12584 15088
rect 13728 15036 13780 15088
rect 13820 15036 13872 15088
rect 14372 15036 14424 15088
rect 17132 15079 17184 15088
rect 17132 15045 17141 15079
rect 17141 15045 17175 15079
rect 17175 15045 17184 15079
rect 17132 15036 17184 15045
rect 17592 15036 17644 15088
rect 12532 14943 12584 14952
rect 12532 14909 12541 14943
rect 12541 14909 12575 14943
rect 12575 14909 12584 14943
rect 12532 14900 12584 14909
rect 12624 14943 12676 14952
rect 12624 14909 12633 14943
rect 12633 14909 12667 14943
rect 12667 14909 12676 14943
rect 12624 14900 12676 14909
rect 12808 14900 12860 14952
rect 12992 14943 13044 14952
rect 12992 14909 13001 14943
rect 13001 14909 13035 14943
rect 13035 14909 13044 14943
rect 12992 14900 13044 14909
rect 15752 14968 15804 15020
rect 13728 14900 13780 14952
rect 13912 14943 13964 14952
rect 13912 14909 13921 14943
rect 13921 14909 13955 14943
rect 13955 14909 13964 14943
rect 13912 14900 13964 14909
rect 14464 14900 14516 14952
rect 15200 14943 15252 14952
rect 15200 14909 15209 14943
rect 15209 14909 15243 14943
rect 15243 14909 15252 14943
rect 15200 14900 15252 14909
rect 15384 14943 15436 14952
rect 15384 14909 15393 14943
rect 15393 14909 15427 14943
rect 15427 14909 15436 14943
rect 15384 14900 15436 14909
rect 15476 14900 15528 14952
rect 16856 14943 16908 14952
rect 16856 14909 16865 14943
rect 16865 14909 16899 14943
rect 16899 14909 16908 14943
rect 16856 14900 16908 14909
rect 17684 14900 17736 14952
rect 12992 14764 13044 14816
rect 13820 14764 13872 14816
rect 14004 14764 14056 14816
rect 14924 14807 14976 14816
rect 14924 14773 14933 14807
rect 14933 14773 14967 14807
rect 14967 14773 14976 14807
rect 14924 14764 14976 14773
rect 15200 14764 15252 14816
rect 15568 14764 15620 14816
rect 15844 14764 15896 14816
rect 17224 14832 17276 14884
rect 17316 14832 17368 14884
rect 16948 14807 17000 14816
rect 16948 14773 16957 14807
rect 16957 14773 16991 14807
rect 16991 14773 17000 14807
rect 16948 14764 17000 14773
rect 4322 14662 4374 14714
rect 4386 14662 4438 14714
rect 4450 14662 4502 14714
rect 4514 14662 4566 14714
rect 4578 14662 4630 14714
rect 12096 14662 12148 14714
rect 12160 14662 12212 14714
rect 12224 14662 12276 14714
rect 12288 14662 12340 14714
rect 12352 14662 12404 14714
rect 19870 14662 19922 14714
rect 19934 14662 19986 14714
rect 19998 14662 20050 14714
rect 20062 14662 20114 14714
rect 20126 14662 20178 14714
rect 27644 14662 27696 14714
rect 27708 14662 27760 14714
rect 27772 14662 27824 14714
rect 27836 14662 27888 14714
rect 27900 14662 27952 14714
rect 14464 14603 14516 14612
rect 14464 14569 14473 14603
rect 14473 14569 14507 14603
rect 14507 14569 14516 14603
rect 14464 14560 14516 14569
rect 14924 14560 14976 14612
rect 12992 14535 13044 14544
rect 12992 14501 13001 14535
rect 13001 14501 13035 14535
rect 13035 14501 13044 14535
rect 12992 14492 13044 14501
rect 13636 14492 13688 14544
rect 14556 14535 14608 14544
rect 14556 14501 14565 14535
rect 14565 14501 14599 14535
rect 14599 14501 14608 14535
rect 17500 14560 17552 14612
rect 18052 14560 18104 14612
rect 18328 14560 18380 14612
rect 14556 14492 14608 14501
rect 12716 14467 12768 14476
rect 12716 14433 12725 14467
rect 12725 14433 12759 14467
rect 12759 14433 12768 14467
rect 12716 14424 12768 14433
rect 13728 14356 13780 14408
rect 15292 14356 15344 14408
rect 16488 14399 16540 14408
rect 16488 14365 16497 14399
rect 16497 14365 16531 14399
rect 16531 14365 16540 14399
rect 16488 14356 16540 14365
rect 16856 14356 16908 14408
rect 17132 14356 17184 14408
rect 17776 14356 17828 14408
rect 14004 14288 14056 14340
rect 31024 14331 31076 14340
rect 31024 14297 31033 14331
rect 31033 14297 31067 14331
rect 31067 14297 31076 14331
rect 31024 14288 31076 14297
rect 15016 14220 15068 14272
rect 3662 14118 3714 14170
rect 3726 14118 3778 14170
rect 3790 14118 3842 14170
rect 3854 14118 3906 14170
rect 3918 14118 3970 14170
rect 11436 14118 11488 14170
rect 11500 14118 11552 14170
rect 11564 14118 11616 14170
rect 11628 14118 11680 14170
rect 11692 14118 11744 14170
rect 19210 14118 19262 14170
rect 19274 14118 19326 14170
rect 19338 14118 19390 14170
rect 19402 14118 19454 14170
rect 19466 14118 19518 14170
rect 26984 14118 27036 14170
rect 27048 14118 27100 14170
rect 27112 14118 27164 14170
rect 27176 14118 27228 14170
rect 27240 14118 27292 14170
rect 13912 14016 13964 14068
rect 16856 14016 16908 14068
rect 16948 14059 17000 14068
rect 16948 14025 16957 14059
rect 16957 14025 16991 14059
rect 16991 14025 17000 14059
rect 16948 14016 17000 14025
rect 13820 13880 13872 13932
rect 15016 13923 15068 13932
rect 15016 13889 15025 13923
rect 15025 13889 15059 13923
rect 15059 13889 15068 13923
rect 15016 13880 15068 13889
rect 15292 13923 15344 13932
rect 15292 13889 15301 13923
rect 15301 13889 15335 13923
rect 15335 13889 15344 13923
rect 15292 13880 15344 13889
rect 18052 13880 18104 13932
rect 17684 13812 17736 13864
rect 17500 13744 17552 13796
rect 4322 13574 4374 13626
rect 4386 13574 4438 13626
rect 4450 13574 4502 13626
rect 4514 13574 4566 13626
rect 4578 13574 4630 13626
rect 12096 13574 12148 13626
rect 12160 13574 12212 13626
rect 12224 13574 12276 13626
rect 12288 13574 12340 13626
rect 12352 13574 12404 13626
rect 19870 13574 19922 13626
rect 19934 13574 19986 13626
rect 19998 13574 20050 13626
rect 20062 13574 20114 13626
rect 20126 13574 20178 13626
rect 27644 13574 27696 13626
rect 27708 13574 27760 13626
rect 27772 13574 27824 13626
rect 27836 13574 27888 13626
rect 27900 13574 27952 13626
rect 3662 13030 3714 13082
rect 3726 13030 3778 13082
rect 3790 13030 3842 13082
rect 3854 13030 3906 13082
rect 3918 13030 3970 13082
rect 11436 13030 11488 13082
rect 11500 13030 11552 13082
rect 11564 13030 11616 13082
rect 11628 13030 11680 13082
rect 11692 13030 11744 13082
rect 19210 13030 19262 13082
rect 19274 13030 19326 13082
rect 19338 13030 19390 13082
rect 19402 13030 19454 13082
rect 19466 13030 19518 13082
rect 26984 13030 27036 13082
rect 27048 13030 27100 13082
rect 27112 13030 27164 13082
rect 27176 13030 27228 13082
rect 27240 13030 27292 13082
rect 4322 12486 4374 12538
rect 4386 12486 4438 12538
rect 4450 12486 4502 12538
rect 4514 12486 4566 12538
rect 4578 12486 4630 12538
rect 12096 12486 12148 12538
rect 12160 12486 12212 12538
rect 12224 12486 12276 12538
rect 12288 12486 12340 12538
rect 12352 12486 12404 12538
rect 19870 12486 19922 12538
rect 19934 12486 19986 12538
rect 19998 12486 20050 12538
rect 20062 12486 20114 12538
rect 20126 12486 20178 12538
rect 27644 12486 27696 12538
rect 27708 12486 27760 12538
rect 27772 12486 27824 12538
rect 27836 12486 27888 12538
rect 27900 12486 27952 12538
rect 3662 11942 3714 11994
rect 3726 11942 3778 11994
rect 3790 11942 3842 11994
rect 3854 11942 3906 11994
rect 3918 11942 3970 11994
rect 11436 11942 11488 11994
rect 11500 11942 11552 11994
rect 11564 11942 11616 11994
rect 11628 11942 11680 11994
rect 11692 11942 11744 11994
rect 19210 11942 19262 11994
rect 19274 11942 19326 11994
rect 19338 11942 19390 11994
rect 19402 11942 19454 11994
rect 19466 11942 19518 11994
rect 26984 11942 27036 11994
rect 27048 11942 27100 11994
rect 27112 11942 27164 11994
rect 27176 11942 27228 11994
rect 27240 11942 27292 11994
rect 4322 11398 4374 11450
rect 4386 11398 4438 11450
rect 4450 11398 4502 11450
rect 4514 11398 4566 11450
rect 4578 11398 4630 11450
rect 12096 11398 12148 11450
rect 12160 11398 12212 11450
rect 12224 11398 12276 11450
rect 12288 11398 12340 11450
rect 12352 11398 12404 11450
rect 19870 11398 19922 11450
rect 19934 11398 19986 11450
rect 19998 11398 20050 11450
rect 20062 11398 20114 11450
rect 20126 11398 20178 11450
rect 27644 11398 27696 11450
rect 27708 11398 27760 11450
rect 27772 11398 27824 11450
rect 27836 11398 27888 11450
rect 27900 11398 27952 11450
rect 3662 10854 3714 10906
rect 3726 10854 3778 10906
rect 3790 10854 3842 10906
rect 3854 10854 3906 10906
rect 3918 10854 3970 10906
rect 11436 10854 11488 10906
rect 11500 10854 11552 10906
rect 11564 10854 11616 10906
rect 11628 10854 11680 10906
rect 11692 10854 11744 10906
rect 19210 10854 19262 10906
rect 19274 10854 19326 10906
rect 19338 10854 19390 10906
rect 19402 10854 19454 10906
rect 19466 10854 19518 10906
rect 26984 10854 27036 10906
rect 27048 10854 27100 10906
rect 27112 10854 27164 10906
rect 27176 10854 27228 10906
rect 27240 10854 27292 10906
rect 4322 10310 4374 10362
rect 4386 10310 4438 10362
rect 4450 10310 4502 10362
rect 4514 10310 4566 10362
rect 4578 10310 4630 10362
rect 12096 10310 12148 10362
rect 12160 10310 12212 10362
rect 12224 10310 12276 10362
rect 12288 10310 12340 10362
rect 12352 10310 12404 10362
rect 19870 10310 19922 10362
rect 19934 10310 19986 10362
rect 19998 10310 20050 10362
rect 20062 10310 20114 10362
rect 20126 10310 20178 10362
rect 27644 10310 27696 10362
rect 27708 10310 27760 10362
rect 27772 10310 27824 10362
rect 27836 10310 27888 10362
rect 27900 10310 27952 10362
rect 3662 9766 3714 9818
rect 3726 9766 3778 9818
rect 3790 9766 3842 9818
rect 3854 9766 3906 9818
rect 3918 9766 3970 9818
rect 11436 9766 11488 9818
rect 11500 9766 11552 9818
rect 11564 9766 11616 9818
rect 11628 9766 11680 9818
rect 11692 9766 11744 9818
rect 19210 9766 19262 9818
rect 19274 9766 19326 9818
rect 19338 9766 19390 9818
rect 19402 9766 19454 9818
rect 19466 9766 19518 9818
rect 26984 9766 27036 9818
rect 27048 9766 27100 9818
rect 27112 9766 27164 9818
rect 27176 9766 27228 9818
rect 27240 9766 27292 9818
rect 4322 9222 4374 9274
rect 4386 9222 4438 9274
rect 4450 9222 4502 9274
rect 4514 9222 4566 9274
rect 4578 9222 4630 9274
rect 12096 9222 12148 9274
rect 12160 9222 12212 9274
rect 12224 9222 12276 9274
rect 12288 9222 12340 9274
rect 12352 9222 12404 9274
rect 19870 9222 19922 9274
rect 19934 9222 19986 9274
rect 19998 9222 20050 9274
rect 20062 9222 20114 9274
rect 20126 9222 20178 9274
rect 27644 9222 27696 9274
rect 27708 9222 27760 9274
rect 27772 9222 27824 9274
rect 27836 9222 27888 9274
rect 27900 9222 27952 9274
rect 3662 8678 3714 8730
rect 3726 8678 3778 8730
rect 3790 8678 3842 8730
rect 3854 8678 3906 8730
rect 3918 8678 3970 8730
rect 11436 8678 11488 8730
rect 11500 8678 11552 8730
rect 11564 8678 11616 8730
rect 11628 8678 11680 8730
rect 11692 8678 11744 8730
rect 19210 8678 19262 8730
rect 19274 8678 19326 8730
rect 19338 8678 19390 8730
rect 19402 8678 19454 8730
rect 19466 8678 19518 8730
rect 26984 8678 27036 8730
rect 27048 8678 27100 8730
rect 27112 8678 27164 8730
rect 27176 8678 27228 8730
rect 27240 8678 27292 8730
rect 4322 8134 4374 8186
rect 4386 8134 4438 8186
rect 4450 8134 4502 8186
rect 4514 8134 4566 8186
rect 4578 8134 4630 8186
rect 12096 8134 12148 8186
rect 12160 8134 12212 8186
rect 12224 8134 12276 8186
rect 12288 8134 12340 8186
rect 12352 8134 12404 8186
rect 19870 8134 19922 8186
rect 19934 8134 19986 8186
rect 19998 8134 20050 8186
rect 20062 8134 20114 8186
rect 20126 8134 20178 8186
rect 27644 8134 27696 8186
rect 27708 8134 27760 8186
rect 27772 8134 27824 8186
rect 27836 8134 27888 8186
rect 27900 8134 27952 8186
rect 3662 7590 3714 7642
rect 3726 7590 3778 7642
rect 3790 7590 3842 7642
rect 3854 7590 3906 7642
rect 3918 7590 3970 7642
rect 11436 7590 11488 7642
rect 11500 7590 11552 7642
rect 11564 7590 11616 7642
rect 11628 7590 11680 7642
rect 11692 7590 11744 7642
rect 19210 7590 19262 7642
rect 19274 7590 19326 7642
rect 19338 7590 19390 7642
rect 19402 7590 19454 7642
rect 19466 7590 19518 7642
rect 26984 7590 27036 7642
rect 27048 7590 27100 7642
rect 27112 7590 27164 7642
rect 27176 7590 27228 7642
rect 27240 7590 27292 7642
rect 4322 7046 4374 7098
rect 4386 7046 4438 7098
rect 4450 7046 4502 7098
rect 4514 7046 4566 7098
rect 4578 7046 4630 7098
rect 12096 7046 12148 7098
rect 12160 7046 12212 7098
rect 12224 7046 12276 7098
rect 12288 7046 12340 7098
rect 12352 7046 12404 7098
rect 19870 7046 19922 7098
rect 19934 7046 19986 7098
rect 19998 7046 20050 7098
rect 20062 7046 20114 7098
rect 20126 7046 20178 7098
rect 27644 7046 27696 7098
rect 27708 7046 27760 7098
rect 27772 7046 27824 7098
rect 27836 7046 27888 7098
rect 27900 7046 27952 7098
rect 3662 6502 3714 6554
rect 3726 6502 3778 6554
rect 3790 6502 3842 6554
rect 3854 6502 3906 6554
rect 3918 6502 3970 6554
rect 11436 6502 11488 6554
rect 11500 6502 11552 6554
rect 11564 6502 11616 6554
rect 11628 6502 11680 6554
rect 11692 6502 11744 6554
rect 19210 6502 19262 6554
rect 19274 6502 19326 6554
rect 19338 6502 19390 6554
rect 19402 6502 19454 6554
rect 19466 6502 19518 6554
rect 26984 6502 27036 6554
rect 27048 6502 27100 6554
rect 27112 6502 27164 6554
rect 27176 6502 27228 6554
rect 27240 6502 27292 6554
rect 4322 5958 4374 6010
rect 4386 5958 4438 6010
rect 4450 5958 4502 6010
rect 4514 5958 4566 6010
rect 4578 5958 4630 6010
rect 12096 5958 12148 6010
rect 12160 5958 12212 6010
rect 12224 5958 12276 6010
rect 12288 5958 12340 6010
rect 12352 5958 12404 6010
rect 19870 5958 19922 6010
rect 19934 5958 19986 6010
rect 19998 5958 20050 6010
rect 20062 5958 20114 6010
rect 20126 5958 20178 6010
rect 27644 5958 27696 6010
rect 27708 5958 27760 6010
rect 27772 5958 27824 6010
rect 27836 5958 27888 6010
rect 27900 5958 27952 6010
rect 3662 5414 3714 5466
rect 3726 5414 3778 5466
rect 3790 5414 3842 5466
rect 3854 5414 3906 5466
rect 3918 5414 3970 5466
rect 11436 5414 11488 5466
rect 11500 5414 11552 5466
rect 11564 5414 11616 5466
rect 11628 5414 11680 5466
rect 11692 5414 11744 5466
rect 19210 5414 19262 5466
rect 19274 5414 19326 5466
rect 19338 5414 19390 5466
rect 19402 5414 19454 5466
rect 19466 5414 19518 5466
rect 26984 5414 27036 5466
rect 27048 5414 27100 5466
rect 27112 5414 27164 5466
rect 27176 5414 27228 5466
rect 27240 5414 27292 5466
rect 4322 4870 4374 4922
rect 4386 4870 4438 4922
rect 4450 4870 4502 4922
rect 4514 4870 4566 4922
rect 4578 4870 4630 4922
rect 12096 4870 12148 4922
rect 12160 4870 12212 4922
rect 12224 4870 12276 4922
rect 12288 4870 12340 4922
rect 12352 4870 12404 4922
rect 19870 4870 19922 4922
rect 19934 4870 19986 4922
rect 19998 4870 20050 4922
rect 20062 4870 20114 4922
rect 20126 4870 20178 4922
rect 27644 4870 27696 4922
rect 27708 4870 27760 4922
rect 27772 4870 27824 4922
rect 27836 4870 27888 4922
rect 27900 4870 27952 4922
rect 3662 4326 3714 4378
rect 3726 4326 3778 4378
rect 3790 4326 3842 4378
rect 3854 4326 3906 4378
rect 3918 4326 3970 4378
rect 11436 4326 11488 4378
rect 11500 4326 11552 4378
rect 11564 4326 11616 4378
rect 11628 4326 11680 4378
rect 11692 4326 11744 4378
rect 19210 4326 19262 4378
rect 19274 4326 19326 4378
rect 19338 4326 19390 4378
rect 19402 4326 19454 4378
rect 19466 4326 19518 4378
rect 26984 4326 27036 4378
rect 27048 4326 27100 4378
rect 27112 4326 27164 4378
rect 27176 4326 27228 4378
rect 27240 4326 27292 4378
rect 4322 3782 4374 3834
rect 4386 3782 4438 3834
rect 4450 3782 4502 3834
rect 4514 3782 4566 3834
rect 4578 3782 4630 3834
rect 12096 3782 12148 3834
rect 12160 3782 12212 3834
rect 12224 3782 12276 3834
rect 12288 3782 12340 3834
rect 12352 3782 12404 3834
rect 19870 3782 19922 3834
rect 19934 3782 19986 3834
rect 19998 3782 20050 3834
rect 20062 3782 20114 3834
rect 20126 3782 20178 3834
rect 27644 3782 27696 3834
rect 27708 3782 27760 3834
rect 27772 3782 27824 3834
rect 27836 3782 27888 3834
rect 27900 3782 27952 3834
rect 3662 3238 3714 3290
rect 3726 3238 3778 3290
rect 3790 3238 3842 3290
rect 3854 3238 3906 3290
rect 3918 3238 3970 3290
rect 11436 3238 11488 3290
rect 11500 3238 11552 3290
rect 11564 3238 11616 3290
rect 11628 3238 11680 3290
rect 11692 3238 11744 3290
rect 19210 3238 19262 3290
rect 19274 3238 19326 3290
rect 19338 3238 19390 3290
rect 19402 3238 19454 3290
rect 19466 3238 19518 3290
rect 26984 3238 27036 3290
rect 27048 3238 27100 3290
rect 27112 3238 27164 3290
rect 27176 3238 27228 3290
rect 27240 3238 27292 3290
rect 4322 2694 4374 2746
rect 4386 2694 4438 2746
rect 4450 2694 4502 2746
rect 4514 2694 4566 2746
rect 4578 2694 4630 2746
rect 12096 2694 12148 2746
rect 12160 2694 12212 2746
rect 12224 2694 12276 2746
rect 12288 2694 12340 2746
rect 12352 2694 12404 2746
rect 19870 2694 19922 2746
rect 19934 2694 19986 2746
rect 19998 2694 20050 2746
rect 20062 2694 20114 2746
rect 20126 2694 20178 2746
rect 27644 2694 27696 2746
rect 27708 2694 27760 2746
rect 27772 2694 27824 2746
rect 27836 2694 27888 2746
rect 27900 2694 27952 2746
rect 3662 2150 3714 2202
rect 3726 2150 3778 2202
rect 3790 2150 3842 2202
rect 3854 2150 3906 2202
rect 3918 2150 3970 2202
rect 11436 2150 11488 2202
rect 11500 2150 11552 2202
rect 11564 2150 11616 2202
rect 11628 2150 11680 2202
rect 11692 2150 11744 2202
rect 19210 2150 19262 2202
rect 19274 2150 19326 2202
rect 19338 2150 19390 2202
rect 19402 2150 19454 2202
rect 19466 2150 19518 2202
rect 26984 2150 27036 2202
rect 27048 2150 27100 2202
rect 27112 2150 27164 2202
rect 27176 2150 27228 2202
rect 27240 2150 27292 2202
rect 4322 1606 4374 1658
rect 4386 1606 4438 1658
rect 4450 1606 4502 1658
rect 4514 1606 4566 1658
rect 4578 1606 4630 1658
rect 12096 1606 12148 1658
rect 12160 1606 12212 1658
rect 12224 1606 12276 1658
rect 12288 1606 12340 1658
rect 12352 1606 12404 1658
rect 19870 1606 19922 1658
rect 19934 1606 19986 1658
rect 19998 1606 20050 1658
rect 20062 1606 20114 1658
rect 20126 1606 20178 1658
rect 27644 1606 27696 1658
rect 27708 1606 27760 1658
rect 27772 1606 27824 1658
rect 27836 1606 27888 1658
rect 27900 1606 27952 1658
rect 3662 1062 3714 1114
rect 3726 1062 3778 1114
rect 3790 1062 3842 1114
rect 3854 1062 3906 1114
rect 3918 1062 3970 1114
rect 11436 1062 11488 1114
rect 11500 1062 11552 1114
rect 11564 1062 11616 1114
rect 11628 1062 11680 1114
rect 11692 1062 11744 1114
rect 19210 1062 19262 1114
rect 19274 1062 19326 1114
rect 19338 1062 19390 1114
rect 19402 1062 19454 1114
rect 19466 1062 19518 1114
rect 26984 1062 27036 1114
rect 27048 1062 27100 1114
rect 27112 1062 27164 1114
rect 27176 1062 27228 1114
rect 27240 1062 27292 1114
rect 17040 1003 17092 1012
rect 17040 969 17049 1003
rect 17049 969 17083 1003
rect 17083 969 17092 1003
rect 17040 960 17092 969
rect 16120 892 16172 944
rect 16764 892 16816 944
rect 7104 756 7156 808
rect 9036 756 9088 808
rect 11612 756 11664 808
rect 12440 756 12492 808
rect 12900 756 12952 808
rect 13544 756 13596 808
rect 14188 756 14240 808
rect 14832 756 14884 808
rect 15476 756 15528 808
rect 16764 756 16816 808
rect 17408 756 17460 808
rect 18052 756 18104 808
rect 18696 756 18748 808
rect 19800 756 19852 808
rect 4322 518 4374 570
rect 4386 518 4438 570
rect 4450 518 4502 570
rect 4514 518 4566 570
rect 4578 518 4630 570
rect 12096 518 12148 570
rect 12160 518 12212 570
rect 12224 518 12276 570
rect 12288 518 12340 570
rect 12352 518 12404 570
rect 19870 518 19922 570
rect 19934 518 19986 570
rect 19998 518 20050 570
rect 20062 518 20114 570
rect 20126 518 20178 570
rect 27644 518 27696 570
rect 27708 518 27760 570
rect 27772 518 27824 570
rect 27836 518 27888 570
rect 27900 518 27952 570
rect 12164 416 12216 468
rect 12440 416 12492 468
<< metal2 >>
rect 10322 19600 10378 20000
rect 11992 19638 12204 19666
rect 4322 19068 4630 19077
rect 4322 19066 4328 19068
rect 4384 19066 4408 19068
rect 4464 19066 4488 19068
rect 4544 19066 4568 19068
rect 4624 19066 4630 19068
rect 4384 19014 4386 19066
rect 4566 19014 4568 19066
rect 4322 19012 4328 19014
rect 4384 19012 4408 19014
rect 4464 19012 4488 19014
rect 4544 19012 4568 19014
rect 4624 19012 4630 19014
rect 4322 19003 4630 19012
rect 10336 18834 10364 19600
rect 11992 18834 12020 19638
rect 12176 19530 12204 19638
rect 12254 19600 12310 20000
rect 12898 19600 12954 20000
rect 13542 19600 13598 20000
rect 14186 19600 14242 20000
rect 14830 19600 14886 20000
rect 16118 19600 16174 20000
rect 16762 19600 16818 20000
rect 17406 19600 17462 20000
rect 22558 19600 22614 20000
rect 12268 19530 12296 19600
rect 12176 19502 12296 19530
rect 12096 19068 12404 19077
rect 12096 19066 12102 19068
rect 12158 19066 12182 19068
rect 12238 19066 12262 19068
rect 12318 19066 12342 19068
rect 12398 19066 12404 19068
rect 12158 19014 12160 19066
rect 12340 19014 12342 19066
rect 12096 19012 12102 19014
rect 12158 19012 12182 19014
rect 12238 19012 12262 19014
rect 12318 19012 12342 19014
rect 12398 19012 12404 19014
rect 12096 19003 12404 19012
rect 12912 18834 12940 19600
rect 13556 18834 13584 19600
rect 14200 18834 14228 19600
rect 14844 18970 14872 19600
rect 16132 18970 16160 19600
rect 14832 18964 14884 18970
rect 14832 18906 14884 18912
rect 16120 18964 16172 18970
rect 16120 18906 16172 18912
rect 10324 18828 10376 18834
rect 10324 18770 10376 18776
rect 11980 18828 12032 18834
rect 11980 18770 12032 18776
rect 12900 18828 12952 18834
rect 12900 18770 12952 18776
rect 13544 18828 13596 18834
rect 13544 18770 13596 18776
rect 14188 18828 14240 18834
rect 14188 18770 14240 18776
rect 15292 18760 15344 18766
rect 15292 18702 15344 18708
rect 848 18624 900 18630
rect 848 18566 900 18572
rect 14372 18624 14424 18630
rect 14372 18566 14424 18572
rect 15200 18624 15252 18630
rect 15200 18566 15252 18572
rect 860 18465 888 18566
rect 3662 18524 3970 18533
rect 3662 18522 3668 18524
rect 3724 18522 3748 18524
rect 3804 18522 3828 18524
rect 3884 18522 3908 18524
rect 3964 18522 3970 18524
rect 3724 18470 3726 18522
rect 3906 18470 3908 18522
rect 3662 18468 3668 18470
rect 3724 18468 3748 18470
rect 3804 18468 3828 18470
rect 3884 18468 3908 18470
rect 3964 18468 3970 18470
rect 846 18456 902 18465
rect 3662 18459 3970 18468
rect 11436 18524 11744 18533
rect 11436 18522 11442 18524
rect 11498 18522 11522 18524
rect 11578 18522 11602 18524
rect 11658 18522 11682 18524
rect 11738 18522 11744 18524
rect 11498 18470 11500 18522
rect 11680 18470 11682 18522
rect 11436 18468 11442 18470
rect 11498 18468 11522 18470
rect 11578 18468 11602 18470
rect 11658 18468 11682 18470
rect 11738 18468 11744 18470
rect 11436 18459 11744 18468
rect 846 18391 902 18400
rect 14188 18284 14240 18290
rect 14188 18226 14240 18232
rect 12716 18216 12768 18222
rect 12716 18158 12768 18164
rect 4322 17980 4630 17989
rect 4322 17978 4328 17980
rect 4384 17978 4408 17980
rect 4464 17978 4488 17980
rect 4544 17978 4568 17980
rect 4624 17978 4630 17980
rect 4384 17926 4386 17978
rect 4566 17926 4568 17978
rect 4322 17924 4328 17926
rect 4384 17924 4408 17926
rect 4464 17924 4488 17926
rect 4544 17924 4568 17926
rect 4624 17924 4630 17926
rect 4322 17915 4630 17924
rect 12096 17980 12404 17989
rect 12096 17978 12102 17980
rect 12158 17978 12182 17980
rect 12238 17978 12262 17980
rect 12318 17978 12342 17980
rect 12398 17978 12404 17980
rect 12158 17926 12160 17978
rect 12340 17926 12342 17978
rect 12096 17924 12102 17926
rect 12158 17924 12182 17926
rect 12238 17924 12262 17926
rect 12318 17924 12342 17926
rect 12398 17924 12404 17926
rect 12096 17915 12404 17924
rect 12532 17672 12584 17678
rect 12532 17614 12584 17620
rect 3662 17436 3970 17445
rect 3662 17434 3668 17436
rect 3724 17434 3748 17436
rect 3804 17434 3828 17436
rect 3884 17434 3908 17436
rect 3964 17434 3970 17436
rect 3724 17382 3726 17434
rect 3906 17382 3908 17434
rect 3662 17380 3668 17382
rect 3724 17380 3748 17382
rect 3804 17380 3828 17382
rect 3884 17380 3908 17382
rect 3964 17380 3970 17382
rect 3662 17371 3970 17380
rect 11436 17436 11744 17445
rect 11436 17434 11442 17436
rect 11498 17434 11522 17436
rect 11578 17434 11602 17436
rect 11658 17434 11682 17436
rect 11738 17434 11744 17436
rect 11498 17382 11500 17434
rect 11680 17382 11682 17434
rect 11436 17380 11442 17382
rect 11498 17380 11522 17382
rect 11578 17380 11602 17382
rect 11658 17380 11682 17382
rect 11738 17380 11744 17382
rect 11436 17371 11744 17380
rect 4322 16892 4630 16901
rect 4322 16890 4328 16892
rect 4384 16890 4408 16892
rect 4464 16890 4488 16892
rect 4544 16890 4568 16892
rect 4624 16890 4630 16892
rect 4384 16838 4386 16890
rect 4566 16838 4568 16890
rect 4322 16836 4328 16838
rect 4384 16836 4408 16838
rect 4464 16836 4488 16838
rect 4544 16836 4568 16838
rect 4624 16836 4630 16838
rect 4322 16827 4630 16836
rect 12096 16892 12404 16901
rect 12096 16890 12102 16892
rect 12158 16890 12182 16892
rect 12238 16890 12262 16892
rect 12318 16890 12342 16892
rect 12398 16890 12404 16892
rect 12158 16838 12160 16890
rect 12340 16838 12342 16890
rect 12096 16836 12102 16838
rect 12158 16836 12182 16838
rect 12238 16836 12262 16838
rect 12318 16836 12342 16838
rect 12398 16836 12404 16838
rect 12096 16827 12404 16836
rect 12544 16658 12572 17614
rect 12728 17542 12756 18158
rect 13636 18080 13688 18086
rect 13636 18022 13688 18028
rect 13648 17746 13676 18022
rect 13636 17740 13688 17746
rect 13636 17682 13688 17688
rect 12716 17536 12768 17542
rect 12716 17478 12768 17484
rect 12728 17270 12756 17478
rect 12716 17264 12768 17270
rect 12716 17206 12768 17212
rect 12728 17066 12756 17206
rect 13648 17202 13676 17682
rect 14200 17542 14228 18226
rect 14384 17785 14412 18566
rect 15212 17814 15240 18566
rect 15304 18426 15332 18702
rect 16776 18698 16804 19600
rect 17316 18828 17368 18834
rect 17316 18770 17368 18776
rect 16764 18692 16816 18698
rect 16764 18634 16816 18640
rect 15384 18624 15436 18630
rect 15384 18566 15436 18572
rect 15292 18420 15344 18426
rect 15292 18362 15344 18368
rect 14740 17808 14792 17814
rect 14370 17776 14426 17785
rect 15200 17808 15252 17814
rect 15014 17776 15070 17785
rect 14792 17756 14872 17762
rect 14740 17750 14872 17756
rect 14370 17711 14426 17720
rect 14648 17740 14700 17746
rect 14384 17678 14412 17711
rect 14752 17734 14872 17750
rect 14648 17682 14700 17688
rect 14372 17672 14424 17678
rect 14372 17614 14424 17620
rect 14660 17610 14688 17682
rect 14648 17604 14700 17610
rect 14648 17546 14700 17552
rect 14004 17536 14056 17542
rect 14004 17478 14056 17484
rect 14188 17536 14240 17542
rect 14188 17478 14240 17484
rect 13636 17196 13688 17202
rect 13636 17138 13688 17144
rect 12716 17060 12768 17066
rect 12716 17002 12768 17008
rect 12532 16652 12584 16658
rect 12532 16594 12584 16600
rect 12728 16590 12756 17002
rect 12716 16584 12768 16590
rect 12716 16526 12768 16532
rect 3662 16348 3970 16357
rect 3662 16346 3668 16348
rect 3724 16346 3748 16348
rect 3804 16346 3828 16348
rect 3884 16346 3908 16348
rect 3964 16346 3970 16348
rect 3724 16294 3726 16346
rect 3906 16294 3908 16346
rect 3662 16292 3668 16294
rect 3724 16292 3748 16294
rect 3804 16292 3828 16294
rect 3884 16292 3908 16294
rect 3964 16292 3970 16294
rect 3662 16283 3970 16292
rect 11436 16348 11744 16357
rect 11436 16346 11442 16348
rect 11498 16346 11522 16348
rect 11578 16346 11602 16348
rect 11658 16346 11682 16348
rect 11738 16346 11744 16348
rect 11498 16294 11500 16346
rect 11680 16294 11682 16346
rect 11436 16292 11442 16294
rect 11498 16292 11522 16294
rect 11578 16292 11602 16294
rect 11658 16292 11682 16294
rect 11738 16292 11744 16294
rect 11436 16283 11744 16292
rect 12532 15904 12584 15910
rect 12532 15846 12584 15852
rect 4322 15804 4630 15813
rect 4322 15802 4328 15804
rect 4384 15802 4408 15804
rect 4464 15802 4488 15804
rect 4544 15802 4568 15804
rect 4624 15802 4630 15804
rect 4384 15750 4386 15802
rect 4566 15750 4568 15802
rect 4322 15748 4328 15750
rect 4384 15748 4408 15750
rect 4464 15748 4488 15750
rect 4544 15748 4568 15750
rect 4624 15748 4630 15750
rect 4322 15739 4630 15748
rect 12096 15804 12404 15813
rect 12096 15802 12102 15804
rect 12158 15802 12182 15804
rect 12238 15802 12262 15804
rect 12318 15802 12342 15804
rect 12398 15802 12404 15804
rect 12158 15750 12160 15802
rect 12340 15750 12342 15802
rect 12096 15748 12102 15750
rect 12158 15748 12182 15750
rect 12238 15748 12262 15750
rect 12318 15748 12342 15750
rect 12398 15748 12404 15750
rect 12096 15739 12404 15748
rect 12544 15638 12572 15846
rect 12532 15632 12584 15638
rect 12532 15574 12584 15580
rect 12728 15366 12756 16526
rect 12808 16244 12860 16250
rect 12808 16186 12860 16192
rect 12716 15360 12768 15366
rect 12716 15302 12768 15308
rect 3662 15260 3970 15269
rect 3662 15258 3668 15260
rect 3724 15258 3748 15260
rect 3804 15258 3828 15260
rect 3884 15258 3908 15260
rect 3964 15258 3970 15260
rect 3724 15206 3726 15258
rect 3906 15206 3908 15258
rect 3662 15204 3668 15206
rect 3724 15204 3748 15206
rect 3804 15204 3828 15206
rect 3884 15204 3908 15206
rect 3964 15204 3970 15206
rect 3662 15195 3970 15204
rect 11436 15260 11744 15269
rect 11436 15258 11442 15260
rect 11498 15258 11522 15260
rect 11578 15258 11602 15260
rect 11658 15258 11682 15260
rect 11738 15258 11744 15260
rect 11498 15206 11500 15258
rect 11680 15206 11682 15258
rect 11436 15204 11442 15206
rect 11498 15204 11522 15206
rect 11578 15204 11602 15206
rect 11658 15204 11682 15206
rect 11738 15204 11744 15206
rect 11436 15195 11744 15204
rect 12624 15156 12676 15162
rect 12624 15098 12676 15104
rect 12532 15088 12584 15094
rect 12532 15030 12584 15036
rect 12544 14958 12572 15030
rect 12636 14958 12664 15098
rect 12532 14952 12584 14958
rect 12532 14894 12584 14900
rect 12624 14952 12676 14958
rect 12624 14894 12676 14900
rect 4322 14716 4630 14725
rect 4322 14714 4328 14716
rect 4384 14714 4408 14716
rect 4464 14714 4488 14716
rect 4544 14714 4568 14716
rect 4624 14714 4630 14716
rect 4384 14662 4386 14714
rect 4566 14662 4568 14714
rect 4322 14660 4328 14662
rect 4384 14660 4408 14662
rect 4464 14660 4488 14662
rect 4544 14660 4568 14662
rect 4624 14660 4630 14662
rect 4322 14651 4630 14660
rect 12096 14716 12404 14725
rect 12096 14714 12102 14716
rect 12158 14714 12182 14716
rect 12238 14714 12262 14716
rect 12318 14714 12342 14716
rect 12398 14714 12404 14716
rect 12158 14662 12160 14714
rect 12340 14662 12342 14714
rect 12096 14660 12102 14662
rect 12158 14660 12182 14662
rect 12238 14660 12262 14662
rect 12318 14660 12342 14662
rect 12398 14660 12404 14662
rect 12096 14651 12404 14660
rect 12728 14482 12756 15302
rect 12820 14958 12848 16186
rect 12992 16040 13044 16046
rect 12992 15982 13044 15988
rect 13004 15502 13032 15982
rect 13648 15570 13676 17138
rect 14016 17134 14044 17478
rect 14660 17338 14688 17546
rect 14648 17332 14700 17338
rect 14648 17274 14700 17280
rect 13728 17128 13780 17134
rect 13728 17070 13780 17076
rect 14004 17128 14056 17134
rect 14004 17070 14056 17076
rect 13740 16046 13768 17070
rect 13820 16992 13872 16998
rect 13820 16934 13872 16940
rect 13832 16046 13860 16934
rect 14016 16522 14044 17070
rect 14844 16998 14872 17734
rect 15200 17750 15252 17756
rect 15014 17711 15016 17720
rect 15068 17711 15070 17720
rect 15016 17682 15068 17688
rect 15292 17672 15344 17678
rect 15292 17614 15344 17620
rect 15108 17332 15160 17338
rect 15108 17274 15160 17280
rect 15120 17218 15148 17274
rect 15120 17190 15240 17218
rect 15304 17202 15332 17614
rect 14188 16992 14240 16998
rect 14188 16934 14240 16940
rect 14832 16992 14884 16998
rect 14832 16934 14884 16940
rect 14200 16794 14228 16934
rect 14188 16788 14240 16794
rect 14188 16730 14240 16736
rect 14844 16658 14872 16934
rect 15212 16658 15240 17190
rect 15292 17196 15344 17202
rect 15292 17138 15344 17144
rect 15396 17066 15424 18566
rect 17328 18426 17356 18770
rect 17420 18442 17448 19600
rect 19870 19068 20178 19077
rect 19870 19066 19876 19068
rect 19932 19066 19956 19068
rect 20012 19066 20036 19068
rect 20092 19066 20116 19068
rect 20172 19066 20178 19068
rect 19932 19014 19934 19066
rect 20114 19014 20116 19066
rect 19870 19012 19876 19014
rect 19932 19012 19956 19014
rect 20012 19012 20036 19014
rect 20092 19012 20116 19014
rect 20172 19012 20178 19014
rect 19870 19003 20178 19012
rect 22572 18834 22600 19600
rect 27644 19068 27952 19077
rect 27644 19066 27650 19068
rect 27706 19066 27730 19068
rect 27786 19066 27810 19068
rect 27866 19066 27890 19068
rect 27946 19066 27952 19068
rect 27706 19014 27708 19066
rect 27888 19014 27890 19066
rect 27644 19012 27650 19014
rect 27706 19012 27730 19014
rect 27786 19012 27810 19014
rect 27866 19012 27890 19014
rect 27946 19012 27952 19014
rect 27644 19003 27952 19012
rect 22560 18828 22612 18834
rect 22560 18770 22612 18776
rect 18236 18624 18288 18630
rect 18236 18566 18288 18572
rect 17420 18426 17540 18442
rect 17316 18420 17368 18426
rect 17420 18420 17552 18426
rect 17420 18414 17500 18420
rect 17316 18362 17368 18368
rect 17500 18362 17552 18368
rect 16396 18284 16448 18290
rect 16396 18226 16448 18232
rect 17132 18284 17184 18290
rect 17132 18226 17184 18232
rect 15844 18216 15896 18222
rect 15844 18158 15896 18164
rect 15856 17882 15884 18158
rect 15844 17876 15896 17882
rect 15844 17818 15896 17824
rect 16304 17672 16356 17678
rect 16304 17614 16356 17620
rect 16316 17338 16344 17614
rect 16304 17332 16356 17338
rect 16304 17274 16356 17280
rect 15384 17060 15436 17066
rect 15384 17002 15436 17008
rect 15476 16788 15528 16794
rect 15476 16730 15528 16736
rect 14832 16652 14884 16658
rect 14832 16594 14884 16600
rect 15200 16652 15252 16658
rect 15200 16594 15252 16600
rect 14004 16516 14056 16522
rect 14004 16458 14056 16464
rect 14016 16182 14044 16458
rect 14556 16244 14608 16250
rect 14556 16186 14608 16192
rect 14004 16176 14056 16182
rect 14056 16124 14136 16130
rect 14004 16118 14136 16124
rect 14016 16102 14136 16118
rect 13728 16040 13780 16046
rect 13728 15982 13780 15988
rect 13820 16040 13872 16046
rect 13820 15982 13872 15988
rect 14004 16040 14056 16046
rect 14004 15982 14056 15988
rect 13636 15564 13688 15570
rect 13636 15506 13688 15512
rect 12992 15496 13044 15502
rect 12992 15438 13044 15444
rect 13004 14958 13032 15438
rect 12808 14952 12860 14958
rect 12808 14894 12860 14900
rect 12992 14952 13044 14958
rect 12992 14894 13044 14900
rect 12992 14816 13044 14822
rect 12992 14758 13044 14764
rect 13004 14550 13032 14758
rect 13648 14550 13676 15506
rect 13740 15450 13768 15982
rect 14016 15706 14044 15982
rect 14108 15706 14136 16102
rect 14372 16108 14424 16114
rect 14372 16050 14424 16056
rect 14384 15978 14412 16050
rect 14372 15972 14424 15978
rect 14372 15914 14424 15920
rect 14004 15700 14056 15706
rect 14004 15642 14056 15648
rect 14096 15700 14148 15706
rect 14096 15642 14148 15648
rect 14384 15570 14412 15914
rect 13820 15564 13872 15570
rect 13820 15506 13872 15512
rect 14372 15564 14424 15570
rect 14372 15506 14424 15512
rect 14464 15564 14516 15570
rect 14464 15506 14516 15512
rect 13832 15450 13860 15506
rect 13740 15422 13860 15450
rect 13912 15428 13964 15434
rect 13740 15094 13768 15422
rect 13912 15370 13964 15376
rect 13728 15088 13780 15094
rect 13728 15030 13780 15036
rect 13820 15088 13872 15094
rect 13820 15030 13872 15036
rect 13740 14958 13768 15030
rect 13728 14952 13780 14958
rect 13728 14894 13780 14900
rect 13832 14822 13860 15030
rect 13924 14958 13952 15370
rect 14384 15094 14412 15506
rect 14372 15088 14424 15094
rect 14372 15030 14424 15036
rect 14476 14958 14504 15506
rect 13912 14952 13964 14958
rect 13912 14894 13964 14900
rect 14464 14952 14516 14958
rect 14464 14894 14516 14900
rect 13820 14816 13872 14822
rect 13820 14758 13872 14764
rect 12992 14544 13044 14550
rect 12992 14486 13044 14492
rect 13636 14544 13688 14550
rect 13688 14492 13860 14498
rect 13636 14486 13860 14492
rect 12716 14476 12768 14482
rect 13648 14470 13860 14486
rect 12716 14418 12768 14424
rect 13740 14414 13768 14470
rect 13728 14408 13780 14414
rect 13728 14350 13780 14356
rect 3662 14172 3970 14181
rect 3662 14170 3668 14172
rect 3724 14170 3748 14172
rect 3804 14170 3828 14172
rect 3884 14170 3908 14172
rect 3964 14170 3970 14172
rect 3724 14118 3726 14170
rect 3906 14118 3908 14170
rect 3662 14116 3668 14118
rect 3724 14116 3748 14118
rect 3804 14116 3828 14118
rect 3884 14116 3908 14118
rect 3964 14116 3970 14118
rect 3662 14107 3970 14116
rect 11436 14172 11744 14181
rect 11436 14170 11442 14172
rect 11498 14170 11522 14172
rect 11578 14170 11602 14172
rect 11658 14170 11682 14172
rect 11738 14170 11744 14172
rect 11498 14118 11500 14170
rect 11680 14118 11682 14170
rect 11436 14116 11442 14118
rect 11498 14116 11522 14118
rect 11578 14116 11602 14118
rect 11658 14116 11682 14118
rect 11738 14116 11744 14118
rect 11436 14107 11744 14116
rect 13832 13938 13860 14470
rect 13924 14074 13952 14894
rect 14004 14816 14056 14822
rect 14004 14758 14056 14764
rect 14016 14346 14044 14758
rect 14476 14618 14504 14894
rect 14464 14612 14516 14618
rect 14464 14554 14516 14560
rect 14568 14550 14596 16186
rect 14740 15700 14792 15706
rect 14740 15642 14792 15648
rect 14752 15366 14780 15642
rect 14924 15564 14976 15570
rect 14924 15506 14976 15512
rect 14936 15434 14964 15506
rect 15212 15434 15240 16594
rect 15488 16250 15516 16730
rect 15568 16652 15620 16658
rect 15568 16594 15620 16600
rect 15580 16522 15608 16594
rect 15568 16516 15620 16522
rect 15568 16458 15620 16464
rect 15844 16448 15896 16454
rect 15844 16390 15896 16396
rect 15476 16244 15528 16250
rect 15476 16186 15528 16192
rect 15752 16108 15804 16114
rect 15752 16050 15804 16056
rect 15764 15570 15792 16050
rect 15856 15638 15884 16390
rect 15844 15632 15896 15638
rect 15844 15574 15896 15580
rect 15476 15564 15528 15570
rect 15476 15506 15528 15512
rect 15752 15564 15804 15570
rect 15752 15506 15804 15512
rect 15936 15564 15988 15570
rect 15936 15506 15988 15512
rect 14924 15428 14976 15434
rect 14924 15370 14976 15376
rect 15200 15428 15252 15434
rect 15200 15370 15252 15376
rect 14740 15360 14792 15366
rect 14740 15302 14792 15308
rect 14752 15162 14780 15302
rect 14740 15156 14792 15162
rect 14740 15098 14792 15104
rect 14936 15042 14964 15370
rect 14936 15014 15424 15042
rect 15396 14958 15424 15014
rect 15488 14958 15516 15506
rect 15568 15496 15620 15502
rect 15568 15438 15620 15444
rect 15200 14952 15252 14958
rect 15200 14894 15252 14900
rect 15384 14952 15436 14958
rect 15384 14894 15436 14900
rect 15476 14952 15528 14958
rect 15476 14894 15528 14900
rect 15212 14822 15240 14894
rect 15580 14822 15608 15438
rect 15764 15026 15792 15506
rect 15948 15162 15976 15506
rect 16408 15450 16436 18226
rect 16764 18216 16816 18222
rect 16764 18158 16816 18164
rect 16776 17542 16804 18158
rect 17144 17746 17172 18226
rect 16856 17740 16908 17746
rect 16856 17682 16908 17688
rect 17132 17740 17184 17746
rect 17132 17682 17184 17688
rect 16764 17536 16816 17542
rect 16764 17478 16816 17484
rect 16776 17338 16804 17478
rect 16868 17338 16896 17682
rect 16764 17332 16816 17338
rect 16764 17274 16816 17280
rect 16856 17332 16908 17338
rect 16856 17274 16908 17280
rect 16672 16992 16724 16998
rect 16672 16934 16724 16940
rect 16684 16726 16712 16934
rect 17144 16726 17172 17682
rect 17328 17678 17356 18362
rect 17684 18080 17736 18086
rect 17684 18022 17736 18028
rect 17776 18080 17828 18086
rect 17776 18022 17828 18028
rect 17316 17672 17368 17678
rect 17316 17614 17368 17620
rect 17592 17672 17644 17678
rect 17592 17614 17644 17620
rect 17408 17536 17460 17542
rect 17408 17478 17460 17484
rect 17420 17066 17448 17478
rect 17604 17338 17632 17614
rect 17592 17332 17644 17338
rect 17592 17274 17644 17280
rect 17696 17218 17724 18022
rect 17788 17338 17816 18022
rect 18248 17882 18276 18566
rect 19210 18524 19518 18533
rect 19210 18522 19216 18524
rect 19272 18522 19296 18524
rect 19352 18522 19376 18524
rect 19432 18522 19456 18524
rect 19512 18522 19518 18524
rect 19272 18470 19274 18522
rect 19454 18470 19456 18522
rect 19210 18468 19216 18470
rect 19272 18468 19296 18470
rect 19352 18468 19376 18470
rect 19432 18468 19456 18470
rect 19512 18468 19518 18470
rect 19210 18459 19518 18468
rect 26984 18524 27292 18533
rect 26984 18522 26990 18524
rect 27046 18522 27070 18524
rect 27126 18522 27150 18524
rect 27206 18522 27230 18524
rect 27286 18522 27292 18524
rect 27046 18470 27048 18522
rect 27228 18470 27230 18522
rect 26984 18468 26990 18470
rect 27046 18468 27070 18470
rect 27126 18468 27150 18470
rect 27206 18468 27230 18470
rect 27286 18468 27292 18470
rect 26984 18459 27292 18468
rect 19870 17980 20178 17989
rect 19870 17978 19876 17980
rect 19932 17978 19956 17980
rect 20012 17978 20036 17980
rect 20092 17978 20116 17980
rect 20172 17978 20178 17980
rect 19932 17926 19934 17978
rect 20114 17926 20116 17978
rect 19870 17924 19876 17926
rect 19932 17924 19956 17926
rect 20012 17924 20036 17926
rect 20092 17924 20116 17926
rect 20172 17924 20178 17926
rect 19870 17915 20178 17924
rect 27644 17980 27952 17989
rect 27644 17978 27650 17980
rect 27706 17978 27730 17980
rect 27786 17978 27810 17980
rect 27866 17978 27890 17980
rect 27946 17978 27952 17980
rect 27706 17926 27708 17978
rect 27888 17926 27890 17978
rect 27644 17924 27650 17926
rect 27706 17924 27730 17926
rect 27786 17924 27810 17926
rect 27866 17924 27890 17926
rect 27946 17924 27952 17926
rect 27644 17915 27952 17924
rect 18236 17876 18288 17882
rect 18236 17818 18288 17824
rect 17960 17808 18012 17814
rect 17960 17750 18012 17756
rect 19064 17808 19116 17814
rect 19064 17750 19116 17756
rect 17776 17332 17828 17338
rect 17776 17274 17828 17280
rect 17696 17190 17908 17218
rect 17316 17060 17368 17066
rect 17316 17002 17368 17008
rect 17408 17060 17460 17066
rect 17408 17002 17460 17008
rect 17684 17060 17736 17066
rect 17684 17002 17736 17008
rect 17328 16726 17356 17002
rect 17500 16992 17552 16998
rect 17500 16934 17552 16940
rect 16672 16720 16724 16726
rect 16672 16662 16724 16668
rect 17132 16720 17184 16726
rect 17132 16662 17184 16668
rect 17316 16720 17368 16726
rect 17316 16662 17368 16668
rect 16580 16652 16632 16658
rect 16500 16612 16580 16640
rect 16500 15570 16528 16612
rect 16580 16594 16632 16600
rect 17040 16652 17092 16658
rect 17040 16594 17092 16600
rect 17224 16652 17276 16658
rect 17224 16594 17276 16600
rect 17052 16538 17080 16594
rect 16948 16516 17000 16522
rect 17052 16510 17172 16538
rect 16948 16458 17000 16464
rect 16672 16448 16724 16454
rect 16672 16390 16724 16396
rect 16684 15570 16712 16390
rect 16764 15972 16816 15978
rect 16764 15914 16816 15920
rect 16488 15564 16540 15570
rect 16488 15506 16540 15512
rect 16672 15564 16724 15570
rect 16672 15506 16724 15512
rect 16408 15434 16528 15450
rect 16408 15428 16540 15434
rect 16408 15422 16488 15428
rect 16488 15370 16540 15376
rect 15936 15156 15988 15162
rect 15936 15098 15988 15104
rect 15752 15020 15804 15026
rect 15752 14962 15804 14968
rect 15948 14906 15976 15098
rect 15856 14878 15976 14906
rect 15856 14822 15884 14878
rect 14924 14816 14976 14822
rect 14924 14758 14976 14764
rect 15200 14816 15252 14822
rect 15200 14758 15252 14764
rect 15568 14816 15620 14822
rect 15568 14758 15620 14764
rect 15844 14816 15896 14822
rect 15844 14758 15896 14764
rect 14936 14618 14964 14758
rect 14924 14612 14976 14618
rect 14924 14554 14976 14560
rect 14556 14544 14608 14550
rect 14556 14486 14608 14492
rect 16500 14414 16528 15370
rect 15292 14408 15344 14414
rect 15292 14350 15344 14356
rect 16488 14408 16540 14414
rect 16488 14350 16540 14356
rect 14004 14340 14056 14346
rect 14004 14282 14056 14288
rect 15016 14272 15068 14278
rect 15016 14214 15068 14220
rect 13912 14068 13964 14074
rect 13912 14010 13964 14016
rect 15028 13938 15056 14214
rect 15304 13938 15332 14350
rect 13820 13932 13872 13938
rect 13820 13874 13872 13880
rect 15016 13932 15068 13938
rect 15016 13874 15068 13880
rect 15292 13932 15344 13938
rect 15292 13874 15344 13880
rect 4322 13628 4630 13637
rect 4322 13626 4328 13628
rect 4384 13626 4408 13628
rect 4464 13626 4488 13628
rect 4544 13626 4568 13628
rect 4624 13626 4630 13628
rect 4384 13574 4386 13626
rect 4566 13574 4568 13626
rect 4322 13572 4328 13574
rect 4384 13572 4408 13574
rect 4464 13572 4488 13574
rect 4544 13572 4568 13574
rect 4624 13572 4630 13574
rect 4322 13563 4630 13572
rect 12096 13628 12404 13637
rect 12096 13626 12102 13628
rect 12158 13626 12182 13628
rect 12238 13626 12262 13628
rect 12318 13626 12342 13628
rect 12398 13626 12404 13628
rect 12158 13574 12160 13626
rect 12340 13574 12342 13626
rect 12096 13572 12102 13574
rect 12158 13572 12182 13574
rect 12238 13572 12262 13574
rect 12318 13572 12342 13574
rect 12398 13572 12404 13574
rect 12096 13563 12404 13572
rect 3662 13084 3970 13093
rect 3662 13082 3668 13084
rect 3724 13082 3748 13084
rect 3804 13082 3828 13084
rect 3884 13082 3908 13084
rect 3964 13082 3970 13084
rect 3724 13030 3726 13082
rect 3906 13030 3908 13082
rect 3662 13028 3668 13030
rect 3724 13028 3748 13030
rect 3804 13028 3828 13030
rect 3884 13028 3908 13030
rect 3964 13028 3970 13030
rect 3662 13019 3970 13028
rect 11436 13084 11744 13093
rect 11436 13082 11442 13084
rect 11498 13082 11522 13084
rect 11578 13082 11602 13084
rect 11658 13082 11682 13084
rect 11738 13082 11744 13084
rect 11498 13030 11500 13082
rect 11680 13030 11682 13082
rect 11436 13028 11442 13030
rect 11498 13028 11522 13030
rect 11578 13028 11602 13030
rect 11658 13028 11682 13030
rect 11738 13028 11744 13030
rect 11436 13019 11744 13028
rect 4322 12540 4630 12549
rect 4322 12538 4328 12540
rect 4384 12538 4408 12540
rect 4464 12538 4488 12540
rect 4544 12538 4568 12540
rect 4624 12538 4630 12540
rect 4384 12486 4386 12538
rect 4566 12486 4568 12538
rect 4322 12484 4328 12486
rect 4384 12484 4408 12486
rect 4464 12484 4488 12486
rect 4544 12484 4568 12486
rect 4624 12484 4630 12486
rect 4322 12475 4630 12484
rect 12096 12540 12404 12549
rect 12096 12538 12102 12540
rect 12158 12538 12182 12540
rect 12238 12538 12262 12540
rect 12318 12538 12342 12540
rect 12398 12538 12404 12540
rect 12158 12486 12160 12538
rect 12340 12486 12342 12538
rect 12096 12484 12102 12486
rect 12158 12484 12182 12486
rect 12238 12484 12262 12486
rect 12318 12484 12342 12486
rect 12398 12484 12404 12486
rect 12096 12475 12404 12484
rect 3662 11996 3970 12005
rect 3662 11994 3668 11996
rect 3724 11994 3748 11996
rect 3804 11994 3828 11996
rect 3884 11994 3908 11996
rect 3964 11994 3970 11996
rect 3724 11942 3726 11994
rect 3906 11942 3908 11994
rect 3662 11940 3668 11942
rect 3724 11940 3748 11942
rect 3804 11940 3828 11942
rect 3884 11940 3908 11942
rect 3964 11940 3970 11942
rect 3662 11931 3970 11940
rect 11436 11996 11744 12005
rect 11436 11994 11442 11996
rect 11498 11994 11522 11996
rect 11578 11994 11602 11996
rect 11658 11994 11682 11996
rect 11738 11994 11744 11996
rect 11498 11942 11500 11994
rect 11680 11942 11682 11994
rect 11436 11940 11442 11942
rect 11498 11940 11522 11942
rect 11578 11940 11602 11942
rect 11658 11940 11682 11942
rect 11738 11940 11744 11942
rect 11436 11931 11744 11940
rect 4322 11452 4630 11461
rect 4322 11450 4328 11452
rect 4384 11450 4408 11452
rect 4464 11450 4488 11452
rect 4544 11450 4568 11452
rect 4624 11450 4630 11452
rect 4384 11398 4386 11450
rect 4566 11398 4568 11450
rect 4322 11396 4328 11398
rect 4384 11396 4408 11398
rect 4464 11396 4488 11398
rect 4544 11396 4568 11398
rect 4624 11396 4630 11398
rect 4322 11387 4630 11396
rect 12096 11452 12404 11461
rect 12096 11450 12102 11452
rect 12158 11450 12182 11452
rect 12238 11450 12262 11452
rect 12318 11450 12342 11452
rect 12398 11450 12404 11452
rect 12158 11398 12160 11450
rect 12340 11398 12342 11450
rect 12096 11396 12102 11398
rect 12158 11396 12182 11398
rect 12238 11396 12262 11398
rect 12318 11396 12342 11398
rect 12398 11396 12404 11398
rect 12096 11387 12404 11396
rect 3662 10908 3970 10917
rect 3662 10906 3668 10908
rect 3724 10906 3748 10908
rect 3804 10906 3828 10908
rect 3884 10906 3908 10908
rect 3964 10906 3970 10908
rect 3724 10854 3726 10906
rect 3906 10854 3908 10906
rect 3662 10852 3668 10854
rect 3724 10852 3748 10854
rect 3804 10852 3828 10854
rect 3884 10852 3908 10854
rect 3964 10852 3970 10854
rect 3662 10843 3970 10852
rect 11436 10908 11744 10917
rect 11436 10906 11442 10908
rect 11498 10906 11522 10908
rect 11578 10906 11602 10908
rect 11658 10906 11682 10908
rect 11738 10906 11744 10908
rect 11498 10854 11500 10906
rect 11680 10854 11682 10906
rect 11436 10852 11442 10854
rect 11498 10852 11522 10854
rect 11578 10852 11602 10854
rect 11658 10852 11682 10854
rect 11738 10852 11744 10854
rect 11436 10843 11744 10852
rect 4322 10364 4630 10373
rect 4322 10362 4328 10364
rect 4384 10362 4408 10364
rect 4464 10362 4488 10364
rect 4544 10362 4568 10364
rect 4624 10362 4630 10364
rect 4384 10310 4386 10362
rect 4566 10310 4568 10362
rect 4322 10308 4328 10310
rect 4384 10308 4408 10310
rect 4464 10308 4488 10310
rect 4544 10308 4568 10310
rect 4624 10308 4630 10310
rect 4322 10299 4630 10308
rect 12096 10364 12404 10373
rect 12096 10362 12102 10364
rect 12158 10362 12182 10364
rect 12238 10362 12262 10364
rect 12318 10362 12342 10364
rect 12398 10362 12404 10364
rect 12158 10310 12160 10362
rect 12340 10310 12342 10362
rect 12096 10308 12102 10310
rect 12158 10308 12182 10310
rect 12238 10308 12262 10310
rect 12318 10308 12342 10310
rect 12398 10308 12404 10310
rect 12096 10299 12404 10308
rect 3662 9820 3970 9829
rect 3662 9818 3668 9820
rect 3724 9818 3748 9820
rect 3804 9818 3828 9820
rect 3884 9818 3908 9820
rect 3964 9818 3970 9820
rect 3724 9766 3726 9818
rect 3906 9766 3908 9818
rect 3662 9764 3668 9766
rect 3724 9764 3748 9766
rect 3804 9764 3828 9766
rect 3884 9764 3908 9766
rect 3964 9764 3970 9766
rect 3662 9755 3970 9764
rect 11436 9820 11744 9829
rect 11436 9818 11442 9820
rect 11498 9818 11522 9820
rect 11578 9818 11602 9820
rect 11658 9818 11682 9820
rect 11738 9818 11744 9820
rect 11498 9766 11500 9818
rect 11680 9766 11682 9818
rect 11436 9764 11442 9766
rect 11498 9764 11522 9766
rect 11578 9764 11602 9766
rect 11658 9764 11682 9766
rect 11738 9764 11744 9766
rect 11436 9755 11744 9764
rect 4322 9276 4630 9285
rect 4322 9274 4328 9276
rect 4384 9274 4408 9276
rect 4464 9274 4488 9276
rect 4544 9274 4568 9276
rect 4624 9274 4630 9276
rect 4384 9222 4386 9274
rect 4566 9222 4568 9274
rect 4322 9220 4328 9222
rect 4384 9220 4408 9222
rect 4464 9220 4488 9222
rect 4544 9220 4568 9222
rect 4624 9220 4630 9222
rect 4322 9211 4630 9220
rect 12096 9276 12404 9285
rect 12096 9274 12102 9276
rect 12158 9274 12182 9276
rect 12238 9274 12262 9276
rect 12318 9274 12342 9276
rect 12398 9274 12404 9276
rect 12158 9222 12160 9274
rect 12340 9222 12342 9274
rect 12096 9220 12102 9222
rect 12158 9220 12182 9222
rect 12238 9220 12262 9222
rect 12318 9220 12342 9222
rect 12398 9220 12404 9222
rect 12096 9211 12404 9220
rect 3662 8732 3970 8741
rect 3662 8730 3668 8732
rect 3724 8730 3748 8732
rect 3804 8730 3828 8732
rect 3884 8730 3908 8732
rect 3964 8730 3970 8732
rect 3724 8678 3726 8730
rect 3906 8678 3908 8730
rect 3662 8676 3668 8678
rect 3724 8676 3748 8678
rect 3804 8676 3828 8678
rect 3884 8676 3908 8678
rect 3964 8676 3970 8678
rect 3662 8667 3970 8676
rect 11436 8732 11744 8741
rect 11436 8730 11442 8732
rect 11498 8730 11522 8732
rect 11578 8730 11602 8732
rect 11658 8730 11682 8732
rect 11738 8730 11744 8732
rect 11498 8678 11500 8730
rect 11680 8678 11682 8730
rect 11436 8676 11442 8678
rect 11498 8676 11522 8678
rect 11578 8676 11602 8678
rect 11658 8676 11682 8678
rect 11738 8676 11744 8678
rect 11436 8667 11744 8676
rect 4322 8188 4630 8197
rect 4322 8186 4328 8188
rect 4384 8186 4408 8188
rect 4464 8186 4488 8188
rect 4544 8186 4568 8188
rect 4624 8186 4630 8188
rect 4384 8134 4386 8186
rect 4566 8134 4568 8186
rect 4322 8132 4328 8134
rect 4384 8132 4408 8134
rect 4464 8132 4488 8134
rect 4544 8132 4568 8134
rect 4624 8132 4630 8134
rect 4322 8123 4630 8132
rect 12096 8188 12404 8197
rect 12096 8186 12102 8188
rect 12158 8186 12182 8188
rect 12238 8186 12262 8188
rect 12318 8186 12342 8188
rect 12398 8186 12404 8188
rect 12158 8134 12160 8186
rect 12340 8134 12342 8186
rect 12096 8132 12102 8134
rect 12158 8132 12182 8134
rect 12238 8132 12262 8134
rect 12318 8132 12342 8134
rect 12398 8132 12404 8134
rect 12096 8123 12404 8132
rect 3662 7644 3970 7653
rect 3662 7642 3668 7644
rect 3724 7642 3748 7644
rect 3804 7642 3828 7644
rect 3884 7642 3908 7644
rect 3964 7642 3970 7644
rect 3724 7590 3726 7642
rect 3906 7590 3908 7642
rect 3662 7588 3668 7590
rect 3724 7588 3748 7590
rect 3804 7588 3828 7590
rect 3884 7588 3908 7590
rect 3964 7588 3970 7590
rect 3662 7579 3970 7588
rect 11436 7644 11744 7653
rect 11436 7642 11442 7644
rect 11498 7642 11522 7644
rect 11578 7642 11602 7644
rect 11658 7642 11682 7644
rect 11738 7642 11744 7644
rect 11498 7590 11500 7642
rect 11680 7590 11682 7642
rect 11436 7588 11442 7590
rect 11498 7588 11522 7590
rect 11578 7588 11602 7590
rect 11658 7588 11682 7590
rect 11738 7588 11744 7590
rect 11436 7579 11744 7588
rect 4322 7100 4630 7109
rect 4322 7098 4328 7100
rect 4384 7098 4408 7100
rect 4464 7098 4488 7100
rect 4544 7098 4568 7100
rect 4624 7098 4630 7100
rect 4384 7046 4386 7098
rect 4566 7046 4568 7098
rect 4322 7044 4328 7046
rect 4384 7044 4408 7046
rect 4464 7044 4488 7046
rect 4544 7044 4568 7046
rect 4624 7044 4630 7046
rect 4322 7035 4630 7044
rect 12096 7100 12404 7109
rect 12096 7098 12102 7100
rect 12158 7098 12182 7100
rect 12238 7098 12262 7100
rect 12318 7098 12342 7100
rect 12398 7098 12404 7100
rect 12158 7046 12160 7098
rect 12340 7046 12342 7098
rect 12096 7044 12102 7046
rect 12158 7044 12182 7046
rect 12238 7044 12262 7046
rect 12318 7044 12342 7046
rect 12398 7044 12404 7046
rect 12096 7035 12404 7044
rect 3662 6556 3970 6565
rect 3662 6554 3668 6556
rect 3724 6554 3748 6556
rect 3804 6554 3828 6556
rect 3884 6554 3908 6556
rect 3964 6554 3970 6556
rect 3724 6502 3726 6554
rect 3906 6502 3908 6554
rect 3662 6500 3668 6502
rect 3724 6500 3748 6502
rect 3804 6500 3828 6502
rect 3884 6500 3908 6502
rect 3964 6500 3970 6502
rect 3662 6491 3970 6500
rect 11436 6556 11744 6565
rect 11436 6554 11442 6556
rect 11498 6554 11522 6556
rect 11578 6554 11602 6556
rect 11658 6554 11682 6556
rect 11738 6554 11744 6556
rect 11498 6502 11500 6554
rect 11680 6502 11682 6554
rect 11436 6500 11442 6502
rect 11498 6500 11522 6502
rect 11578 6500 11602 6502
rect 11658 6500 11682 6502
rect 11738 6500 11744 6502
rect 11436 6491 11744 6500
rect 4322 6012 4630 6021
rect 4322 6010 4328 6012
rect 4384 6010 4408 6012
rect 4464 6010 4488 6012
rect 4544 6010 4568 6012
rect 4624 6010 4630 6012
rect 4384 5958 4386 6010
rect 4566 5958 4568 6010
rect 4322 5956 4328 5958
rect 4384 5956 4408 5958
rect 4464 5956 4488 5958
rect 4544 5956 4568 5958
rect 4624 5956 4630 5958
rect 4322 5947 4630 5956
rect 12096 6012 12404 6021
rect 12096 6010 12102 6012
rect 12158 6010 12182 6012
rect 12238 6010 12262 6012
rect 12318 6010 12342 6012
rect 12398 6010 12404 6012
rect 12158 5958 12160 6010
rect 12340 5958 12342 6010
rect 12096 5956 12102 5958
rect 12158 5956 12182 5958
rect 12238 5956 12262 5958
rect 12318 5956 12342 5958
rect 12398 5956 12404 5958
rect 12096 5947 12404 5956
rect 3662 5468 3970 5477
rect 3662 5466 3668 5468
rect 3724 5466 3748 5468
rect 3804 5466 3828 5468
rect 3884 5466 3908 5468
rect 3964 5466 3970 5468
rect 3724 5414 3726 5466
rect 3906 5414 3908 5466
rect 3662 5412 3668 5414
rect 3724 5412 3748 5414
rect 3804 5412 3828 5414
rect 3884 5412 3908 5414
rect 3964 5412 3970 5414
rect 3662 5403 3970 5412
rect 11436 5468 11744 5477
rect 11436 5466 11442 5468
rect 11498 5466 11522 5468
rect 11578 5466 11602 5468
rect 11658 5466 11682 5468
rect 11738 5466 11744 5468
rect 11498 5414 11500 5466
rect 11680 5414 11682 5466
rect 11436 5412 11442 5414
rect 11498 5412 11522 5414
rect 11578 5412 11602 5414
rect 11658 5412 11682 5414
rect 11738 5412 11744 5414
rect 11436 5403 11744 5412
rect 4322 4924 4630 4933
rect 4322 4922 4328 4924
rect 4384 4922 4408 4924
rect 4464 4922 4488 4924
rect 4544 4922 4568 4924
rect 4624 4922 4630 4924
rect 4384 4870 4386 4922
rect 4566 4870 4568 4922
rect 4322 4868 4328 4870
rect 4384 4868 4408 4870
rect 4464 4868 4488 4870
rect 4544 4868 4568 4870
rect 4624 4868 4630 4870
rect 4322 4859 4630 4868
rect 12096 4924 12404 4933
rect 12096 4922 12102 4924
rect 12158 4922 12182 4924
rect 12238 4922 12262 4924
rect 12318 4922 12342 4924
rect 12398 4922 12404 4924
rect 12158 4870 12160 4922
rect 12340 4870 12342 4922
rect 12096 4868 12102 4870
rect 12158 4868 12182 4870
rect 12238 4868 12262 4870
rect 12318 4868 12342 4870
rect 12398 4868 12404 4870
rect 12096 4859 12404 4868
rect 3662 4380 3970 4389
rect 3662 4378 3668 4380
rect 3724 4378 3748 4380
rect 3804 4378 3828 4380
rect 3884 4378 3908 4380
rect 3964 4378 3970 4380
rect 3724 4326 3726 4378
rect 3906 4326 3908 4378
rect 3662 4324 3668 4326
rect 3724 4324 3748 4326
rect 3804 4324 3828 4326
rect 3884 4324 3908 4326
rect 3964 4324 3970 4326
rect 3662 4315 3970 4324
rect 11436 4380 11744 4389
rect 11436 4378 11442 4380
rect 11498 4378 11522 4380
rect 11578 4378 11602 4380
rect 11658 4378 11682 4380
rect 11738 4378 11744 4380
rect 11498 4326 11500 4378
rect 11680 4326 11682 4378
rect 11436 4324 11442 4326
rect 11498 4324 11522 4326
rect 11578 4324 11602 4326
rect 11658 4324 11682 4326
rect 11738 4324 11744 4326
rect 11436 4315 11744 4324
rect 4322 3836 4630 3845
rect 4322 3834 4328 3836
rect 4384 3834 4408 3836
rect 4464 3834 4488 3836
rect 4544 3834 4568 3836
rect 4624 3834 4630 3836
rect 4384 3782 4386 3834
rect 4566 3782 4568 3834
rect 4322 3780 4328 3782
rect 4384 3780 4408 3782
rect 4464 3780 4488 3782
rect 4544 3780 4568 3782
rect 4624 3780 4630 3782
rect 4322 3771 4630 3780
rect 12096 3836 12404 3845
rect 12096 3834 12102 3836
rect 12158 3834 12182 3836
rect 12238 3834 12262 3836
rect 12318 3834 12342 3836
rect 12398 3834 12404 3836
rect 12158 3782 12160 3834
rect 12340 3782 12342 3834
rect 12096 3780 12102 3782
rect 12158 3780 12182 3782
rect 12238 3780 12262 3782
rect 12318 3780 12342 3782
rect 12398 3780 12404 3782
rect 12096 3771 12404 3780
rect 3662 3292 3970 3301
rect 3662 3290 3668 3292
rect 3724 3290 3748 3292
rect 3804 3290 3828 3292
rect 3884 3290 3908 3292
rect 3964 3290 3970 3292
rect 3724 3238 3726 3290
rect 3906 3238 3908 3290
rect 3662 3236 3668 3238
rect 3724 3236 3748 3238
rect 3804 3236 3828 3238
rect 3884 3236 3908 3238
rect 3964 3236 3970 3238
rect 3662 3227 3970 3236
rect 11436 3292 11744 3301
rect 11436 3290 11442 3292
rect 11498 3290 11522 3292
rect 11578 3290 11602 3292
rect 11658 3290 11682 3292
rect 11738 3290 11744 3292
rect 11498 3238 11500 3290
rect 11680 3238 11682 3290
rect 11436 3236 11442 3238
rect 11498 3236 11522 3238
rect 11578 3236 11602 3238
rect 11658 3236 11682 3238
rect 11738 3236 11744 3238
rect 11436 3227 11744 3236
rect 4322 2748 4630 2757
rect 4322 2746 4328 2748
rect 4384 2746 4408 2748
rect 4464 2746 4488 2748
rect 4544 2746 4568 2748
rect 4624 2746 4630 2748
rect 4384 2694 4386 2746
rect 4566 2694 4568 2746
rect 4322 2692 4328 2694
rect 4384 2692 4408 2694
rect 4464 2692 4488 2694
rect 4544 2692 4568 2694
rect 4624 2692 4630 2694
rect 4322 2683 4630 2692
rect 12096 2748 12404 2757
rect 12096 2746 12102 2748
rect 12158 2746 12182 2748
rect 12238 2746 12262 2748
rect 12318 2746 12342 2748
rect 12398 2746 12404 2748
rect 12158 2694 12160 2746
rect 12340 2694 12342 2746
rect 12096 2692 12102 2694
rect 12158 2692 12182 2694
rect 12238 2692 12262 2694
rect 12318 2692 12342 2694
rect 12398 2692 12404 2694
rect 12096 2683 12404 2692
rect 3662 2204 3970 2213
rect 3662 2202 3668 2204
rect 3724 2202 3748 2204
rect 3804 2202 3828 2204
rect 3884 2202 3908 2204
rect 3964 2202 3970 2204
rect 3724 2150 3726 2202
rect 3906 2150 3908 2202
rect 3662 2148 3668 2150
rect 3724 2148 3748 2150
rect 3804 2148 3828 2150
rect 3884 2148 3908 2150
rect 3964 2148 3970 2150
rect 3662 2139 3970 2148
rect 11436 2204 11744 2213
rect 11436 2202 11442 2204
rect 11498 2202 11522 2204
rect 11578 2202 11602 2204
rect 11658 2202 11682 2204
rect 11738 2202 11744 2204
rect 11498 2150 11500 2202
rect 11680 2150 11682 2202
rect 11436 2148 11442 2150
rect 11498 2148 11522 2150
rect 11578 2148 11602 2150
rect 11658 2148 11682 2150
rect 11738 2148 11744 2150
rect 11436 2139 11744 2148
rect 4322 1660 4630 1669
rect 4322 1658 4328 1660
rect 4384 1658 4408 1660
rect 4464 1658 4488 1660
rect 4544 1658 4568 1660
rect 4624 1658 4630 1660
rect 4384 1606 4386 1658
rect 4566 1606 4568 1658
rect 4322 1604 4328 1606
rect 4384 1604 4408 1606
rect 4464 1604 4488 1606
rect 4544 1604 4568 1606
rect 4624 1604 4630 1606
rect 4322 1595 4630 1604
rect 12096 1660 12404 1669
rect 12096 1658 12102 1660
rect 12158 1658 12182 1660
rect 12238 1658 12262 1660
rect 12318 1658 12342 1660
rect 12398 1658 12404 1660
rect 12158 1606 12160 1658
rect 12340 1606 12342 1658
rect 12096 1604 12102 1606
rect 12158 1604 12182 1606
rect 12238 1604 12262 1606
rect 12318 1604 12342 1606
rect 12398 1604 12404 1606
rect 12096 1595 12404 1604
rect 3662 1116 3970 1125
rect 3662 1114 3668 1116
rect 3724 1114 3748 1116
rect 3804 1114 3828 1116
rect 3884 1114 3908 1116
rect 3964 1114 3970 1116
rect 3724 1062 3726 1114
rect 3906 1062 3908 1114
rect 3662 1060 3668 1062
rect 3724 1060 3748 1062
rect 3804 1060 3828 1062
rect 3884 1060 3908 1062
rect 3964 1060 3970 1062
rect 3662 1051 3970 1060
rect 11436 1116 11744 1125
rect 11436 1114 11442 1116
rect 11498 1114 11522 1116
rect 11578 1114 11602 1116
rect 11658 1114 11682 1116
rect 11738 1114 11744 1116
rect 11498 1062 11500 1114
rect 11680 1062 11682 1114
rect 11436 1060 11442 1062
rect 11498 1060 11522 1062
rect 11578 1060 11602 1062
rect 11658 1060 11682 1062
rect 11738 1060 11744 1062
rect 11436 1051 11744 1060
rect 16776 950 16804 15914
rect 16856 15904 16908 15910
rect 16856 15846 16908 15852
rect 16868 14958 16896 15846
rect 16960 15706 16988 16458
rect 17040 16448 17092 16454
rect 17040 16390 17092 16396
rect 17052 16046 17080 16390
rect 17040 16040 17092 16046
rect 17040 15982 17092 15988
rect 16948 15700 17000 15706
rect 16948 15642 17000 15648
rect 17052 15366 17080 15982
rect 17144 15910 17172 16510
rect 17236 16046 17264 16594
rect 17224 16040 17276 16046
rect 17224 15982 17276 15988
rect 17132 15904 17184 15910
rect 17132 15846 17184 15852
rect 17132 15564 17184 15570
rect 17132 15506 17184 15512
rect 17040 15360 17092 15366
rect 17040 15302 17092 15308
rect 17052 15162 17080 15302
rect 17040 15156 17092 15162
rect 17040 15098 17092 15104
rect 17144 15094 17172 15506
rect 17132 15088 17184 15094
rect 17132 15030 17184 15036
rect 16856 14952 16908 14958
rect 16856 14894 16908 14900
rect 17236 14890 17264 15982
rect 17316 15904 17368 15910
rect 17316 15846 17368 15852
rect 17408 15904 17460 15910
rect 17408 15846 17460 15852
rect 17328 14890 17356 15846
rect 17420 15570 17448 15846
rect 17512 15706 17540 16934
rect 17592 15904 17644 15910
rect 17592 15846 17644 15852
rect 17500 15700 17552 15706
rect 17500 15642 17552 15648
rect 17408 15564 17460 15570
rect 17408 15506 17460 15512
rect 17512 15162 17540 15642
rect 17500 15156 17552 15162
rect 17500 15098 17552 15104
rect 17224 14884 17276 14890
rect 17224 14826 17276 14832
rect 17316 14884 17368 14890
rect 17316 14826 17368 14832
rect 16948 14816 17000 14822
rect 16948 14758 17000 14764
rect 16856 14408 16908 14414
rect 16856 14350 16908 14356
rect 16868 14074 16896 14350
rect 16960 14074 16988 14758
rect 17512 14618 17540 15098
rect 17604 15094 17632 15846
rect 17592 15088 17644 15094
rect 17592 15030 17644 15036
rect 17696 14958 17724 17002
rect 17880 15586 17908 17190
rect 17972 17134 18000 17750
rect 18328 17196 18380 17202
rect 18328 17138 18380 17144
rect 17960 17128 18012 17134
rect 17960 17070 18012 17076
rect 17972 15638 18000 17070
rect 18236 16176 18288 16182
rect 18340 16130 18368 17138
rect 18880 16584 18932 16590
rect 18880 16526 18932 16532
rect 19076 16538 19104 17750
rect 19210 17436 19518 17445
rect 19210 17434 19216 17436
rect 19272 17434 19296 17436
rect 19352 17434 19376 17436
rect 19432 17434 19456 17436
rect 19512 17434 19518 17436
rect 19272 17382 19274 17434
rect 19454 17382 19456 17434
rect 19210 17380 19216 17382
rect 19272 17380 19296 17382
rect 19352 17380 19376 17382
rect 19432 17380 19456 17382
rect 19512 17380 19518 17382
rect 19210 17371 19518 17380
rect 26984 17436 27292 17445
rect 26984 17434 26990 17436
rect 27046 17434 27070 17436
rect 27126 17434 27150 17436
rect 27206 17434 27230 17436
rect 27286 17434 27292 17436
rect 27046 17382 27048 17434
rect 27228 17382 27230 17434
rect 26984 17380 26990 17382
rect 27046 17380 27070 17382
rect 27126 17380 27150 17382
rect 27206 17380 27230 17382
rect 27286 17380 27292 17382
rect 26984 17371 27292 17380
rect 19870 16892 20178 16901
rect 19870 16890 19876 16892
rect 19932 16890 19956 16892
rect 20012 16890 20036 16892
rect 20092 16890 20116 16892
rect 20172 16890 20178 16892
rect 19932 16838 19934 16890
rect 20114 16838 20116 16890
rect 19870 16836 19876 16838
rect 19932 16836 19956 16838
rect 20012 16836 20036 16838
rect 20092 16836 20116 16838
rect 20172 16836 20178 16838
rect 19870 16827 20178 16836
rect 27644 16892 27952 16901
rect 27644 16890 27650 16892
rect 27706 16890 27730 16892
rect 27786 16890 27810 16892
rect 27866 16890 27890 16892
rect 27946 16890 27952 16892
rect 27706 16838 27708 16890
rect 27888 16838 27890 16890
rect 27644 16836 27650 16838
rect 27706 16836 27730 16838
rect 27786 16836 27810 16838
rect 27866 16836 27890 16838
rect 27946 16836 27952 16838
rect 27644 16827 27952 16836
rect 19156 16652 19208 16658
rect 19156 16594 19208 16600
rect 19168 16538 19196 16594
rect 18288 16124 18368 16130
rect 18236 16118 18368 16124
rect 18248 16102 18368 16118
rect 18340 15978 18368 16102
rect 18052 15972 18104 15978
rect 18052 15914 18104 15920
rect 18328 15972 18380 15978
rect 18328 15914 18380 15920
rect 17788 15558 17908 15586
rect 17960 15632 18012 15638
rect 17960 15574 18012 15580
rect 17684 14952 17736 14958
rect 17684 14894 17736 14900
rect 17500 14612 17552 14618
rect 17500 14554 17552 14560
rect 17132 14408 17184 14414
rect 17132 14350 17184 14356
rect 16856 14068 16908 14074
rect 16856 14010 16908 14016
rect 16948 14068 17000 14074
rect 16948 14010 17000 14016
rect 17144 6914 17172 14350
rect 17512 13802 17540 14554
rect 17696 13870 17724 14894
rect 17788 14414 17816 15558
rect 17868 15496 17920 15502
rect 17868 15438 17920 15444
rect 17880 15162 17908 15438
rect 17868 15156 17920 15162
rect 17868 15098 17920 15104
rect 18064 14618 18092 15914
rect 18892 15706 18920 16526
rect 19076 16522 19196 16538
rect 19076 16516 19208 16522
rect 19076 16510 19156 16516
rect 18880 15700 18932 15706
rect 18880 15642 18932 15648
rect 18328 15632 18380 15638
rect 18328 15574 18380 15580
rect 18340 14618 18368 15574
rect 19076 15366 19104 16510
rect 19156 16458 19208 16464
rect 19210 16348 19518 16357
rect 19210 16346 19216 16348
rect 19272 16346 19296 16348
rect 19352 16346 19376 16348
rect 19432 16346 19456 16348
rect 19512 16346 19518 16348
rect 19272 16294 19274 16346
rect 19454 16294 19456 16346
rect 19210 16292 19216 16294
rect 19272 16292 19296 16294
rect 19352 16292 19376 16294
rect 19432 16292 19456 16294
rect 19512 16292 19518 16294
rect 19210 16283 19518 16292
rect 26984 16348 27292 16357
rect 26984 16346 26990 16348
rect 27046 16346 27070 16348
rect 27126 16346 27150 16348
rect 27206 16346 27230 16348
rect 27286 16346 27292 16348
rect 27046 16294 27048 16346
rect 27228 16294 27230 16346
rect 26984 16292 26990 16294
rect 27046 16292 27070 16294
rect 27126 16292 27150 16294
rect 27206 16292 27230 16294
rect 27286 16292 27292 16294
rect 26984 16283 27292 16292
rect 19340 16244 19392 16250
rect 19340 16186 19392 16192
rect 19352 15706 19380 16186
rect 19870 15804 20178 15813
rect 19870 15802 19876 15804
rect 19932 15802 19956 15804
rect 20012 15802 20036 15804
rect 20092 15802 20116 15804
rect 20172 15802 20178 15804
rect 19932 15750 19934 15802
rect 20114 15750 20116 15802
rect 19870 15748 19876 15750
rect 19932 15748 19956 15750
rect 20012 15748 20036 15750
rect 20092 15748 20116 15750
rect 20172 15748 20178 15750
rect 19870 15739 20178 15748
rect 27644 15804 27952 15813
rect 27644 15802 27650 15804
rect 27706 15802 27730 15804
rect 27786 15802 27810 15804
rect 27866 15802 27890 15804
rect 27946 15802 27952 15804
rect 27706 15750 27708 15802
rect 27888 15750 27890 15802
rect 27644 15748 27650 15750
rect 27706 15748 27730 15750
rect 27786 15748 27810 15750
rect 27866 15748 27890 15750
rect 27946 15748 27952 15750
rect 27644 15739 27952 15748
rect 19340 15700 19392 15706
rect 19340 15642 19392 15648
rect 19064 15360 19116 15366
rect 19064 15302 19116 15308
rect 19210 15260 19518 15269
rect 19210 15258 19216 15260
rect 19272 15258 19296 15260
rect 19352 15258 19376 15260
rect 19432 15258 19456 15260
rect 19512 15258 19518 15260
rect 19272 15206 19274 15258
rect 19454 15206 19456 15258
rect 19210 15204 19216 15206
rect 19272 15204 19296 15206
rect 19352 15204 19376 15206
rect 19432 15204 19456 15206
rect 19512 15204 19518 15206
rect 19210 15195 19518 15204
rect 26984 15260 27292 15269
rect 26984 15258 26990 15260
rect 27046 15258 27070 15260
rect 27126 15258 27150 15260
rect 27206 15258 27230 15260
rect 27286 15258 27292 15260
rect 27046 15206 27048 15258
rect 27228 15206 27230 15258
rect 26984 15204 26990 15206
rect 27046 15204 27070 15206
rect 27126 15204 27150 15206
rect 27206 15204 27230 15206
rect 27286 15204 27292 15206
rect 26984 15195 27292 15204
rect 19870 14716 20178 14725
rect 19870 14714 19876 14716
rect 19932 14714 19956 14716
rect 20012 14714 20036 14716
rect 20092 14714 20116 14716
rect 20172 14714 20178 14716
rect 19932 14662 19934 14714
rect 20114 14662 20116 14714
rect 19870 14660 19876 14662
rect 19932 14660 19956 14662
rect 20012 14660 20036 14662
rect 20092 14660 20116 14662
rect 20172 14660 20178 14662
rect 19870 14651 20178 14660
rect 27644 14716 27952 14725
rect 27644 14714 27650 14716
rect 27706 14714 27730 14716
rect 27786 14714 27810 14716
rect 27866 14714 27890 14716
rect 27946 14714 27952 14716
rect 27706 14662 27708 14714
rect 27888 14662 27890 14714
rect 27644 14660 27650 14662
rect 27706 14660 27730 14662
rect 27786 14660 27810 14662
rect 27866 14660 27890 14662
rect 27946 14660 27952 14662
rect 27644 14651 27952 14660
rect 18052 14612 18104 14618
rect 18052 14554 18104 14560
rect 18328 14612 18380 14618
rect 18328 14554 18380 14560
rect 17776 14408 17828 14414
rect 17776 14350 17828 14356
rect 18064 13938 18092 14554
rect 31022 14376 31078 14385
rect 31022 14311 31024 14320
rect 31076 14311 31078 14320
rect 31024 14282 31076 14288
rect 19210 14172 19518 14181
rect 19210 14170 19216 14172
rect 19272 14170 19296 14172
rect 19352 14170 19376 14172
rect 19432 14170 19456 14172
rect 19512 14170 19518 14172
rect 19272 14118 19274 14170
rect 19454 14118 19456 14170
rect 19210 14116 19216 14118
rect 19272 14116 19296 14118
rect 19352 14116 19376 14118
rect 19432 14116 19456 14118
rect 19512 14116 19518 14118
rect 19210 14107 19518 14116
rect 26984 14172 27292 14181
rect 26984 14170 26990 14172
rect 27046 14170 27070 14172
rect 27126 14170 27150 14172
rect 27206 14170 27230 14172
rect 27286 14170 27292 14172
rect 27046 14118 27048 14170
rect 27228 14118 27230 14170
rect 26984 14116 26990 14118
rect 27046 14116 27070 14118
rect 27126 14116 27150 14118
rect 27206 14116 27230 14118
rect 27286 14116 27292 14118
rect 26984 14107 27292 14116
rect 18052 13932 18104 13938
rect 18052 13874 18104 13880
rect 17684 13864 17736 13870
rect 17684 13806 17736 13812
rect 17500 13796 17552 13802
rect 17500 13738 17552 13744
rect 19870 13628 20178 13637
rect 19870 13626 19876 13628
rect 19932 13626 19956 13628
rect 20012 13626 20036 13628
rect 20092 13626 20116 13628
rect 20172 13626 20178 13628
rect 19932 13574 19934 13626
rect 20114 13574 20116 13626
rect 19870 13572 19876 13574
rect 19932 13572 19956 13574
rect 20012 13572 20036 13574
rect 20092 13572 20116 13574
rect 20172 13572 20178 13574
rect 19870 13563 20178 13572
rect 27644 13628 27952 13637
rect 27644 13626 27650 13628
rect 27706 13626 27730 13628
rect 27786 13626 27810 13628
rect 27866 13626 27890 13628
rect 27946 13626 27952 13628
rect 27706 13574 27708 13626
rect 27888 13574 27890 13626
rect 27644 13572 27650 13574
rect 27706 13572 27730 13574
rect 27786 13572 27810 13574
rect 27866 13572 27890 13574
rect 27946 13572 27952 13574
rect 27644 13563 27952 13572
rect 19210 13084 19518 13093
rect 19210 13082 19216 13084
rect 19272 13082 19296 13084
rect 19352 13082 19376 13084
rect 19432 13082 19456 13084
rect 19512 13082 19518 13084
rect 19272 13030 19274 13082
rect 19454 13030 19456 13082
rect 19210 13028 19216 13030
rect 19272 13028 19296 13030
rect 19352 13028 19376 13030
rect 19432 13028 19456 13030
rect 19512 13028 19518 13030
rect 19210 13019 19518 13028
rect 26984 13084 27292 13093
rect 26984 13082 26990 13084
rect 27046 13082 27070 13084
rect 27126 13082 27150 13084
rect 27206 13082 27230 13084
rect 27286 13082 27292 13084
rect 27046 13030 27048 13082
rect 27228 13030 27230 13082
rect 26984 13028 26990 13030
rect 27046 13028 27070 13030
rect 27126 13028 27150 13030
rect 27206 13028 27230 13030
rect 27286 13028 27292 13030
rect 26984 13019 27292 13028
rect 19870 12540 20178 12549
rect 19870 12538 19876 12540
rect 19932 12538 19956 12540
rect 20012 12538 20036 12540
rect 20092 12538 20116 12540
rect 20172 12538 20178 12540
rect 19932 12486 19934 12538
rect 20114 12486 20116 12538
rect 19870 12484 19876 12486
rect 19932 12484 19956 12486
rect 20012 12484 20036 12486
rect 20092 12484 20116 12486
rect 20172 12484 20178 12486
rect 19870 12475 20178 12484
rect 27644 12540 27952 12549
rect 27644 12538 27650 12540
rect 27706 12538 27730 12540
rect 27786 12538 27810 12540
rect 27866 12538 27890 12540
rect 27946 12538 27952 12540
rect 27706 12486 27708 12538
rect 27888 12486 27890 12538
rect 27644 12484 27650 12486
rect 27706 12484 27730 12486
rect 27786 12484 27810 12486
rect 27866 12484 27890 12486
rect 27946 12484 27952 12486
rect 27644 12475 27952 12484
rect 19210 11996 19518 12005
rect 19210 11994 19216 11996
rect 19272 11994 19296 11996
rect 19352 11994 19376 11996
rect 19432 11994 19456 11996
rect 19512 11994 19518 11996
rect 19272 11942 19274 11994
rect 19454 11942 19456 11994
rect 19210 11940 19216 11942
rect 19272 11940 19296 11942
rect 19352 11940 19376 11942
rect 19432 11940 19456 11942
rect 19512 11940 19518 11942
rect 19210 11931 19518 11940
rect 26984 11996 27292 12005
rect 26984 11994 26990 11996
rect 27046 11994 27070 11996
rect 27126 11994 27150 11996
rect 27206 11994 27230 11996
rect 27286 11994 27292 11996
rect 27046 11942 27048 11994
rect 27228 11942 27230 11994
rect 26984 11940 26990 11942
rect 27046 11940 27070 11942
rect 27126 11940 27150 11942
rect 27206 11940 27230 11942
rect 27286 11940 27292 11942
rect 26984 11931 27292 11940
rect 19870 11452 20178 11461
rect 19870 11450 19876 11452
rect 19932 11450 19956 11452
rect 20012 11450 20036 11452
rect 20092 11450 20116 11452
rect 20172 11450 20178 11452
rect 19932 11398 19934 11450
rect 20114 11398 20116 11450
rect 19870 11396 19876 11398
rect 19932 11396 19956 11398
rect 20012 11396 20036 11398
rect 20092 11396 20116 11398
rect 20172 11396 20178 11398
rect 19870 11387 20178 11396
rect 27644 11452 27952 11461
rect 27644 11450 27650 11452
rect 27706 11450 27730 11452
rect 27786 11450 27810 11452
rect 27866 11450 27890 11452
rect 27946 11450 27952 11452
rect 27706 11398 27708 11450
rect 27888 11398 27890 11450
rect 27644 11396 27650 11398
rect 27706 11396 27730 11398
rect 27786 11396 27810 11398
rect 27866 11396 27890 11398
rect 27946 11396 27952 11398
rect 27644 11387 27952 11396
rect 19210 10908 19518 10917
rect 19210 10906 19216 10908
rect 19272 10906 19296 10908
rect 19352 10906 19376 10908
rect 19432 10906 19456 10908
rect 19512 10906 19518 10908
rect 19272 10854 19274 10906
rect 19454 10854 19456 10906
rect 19210 10852 19216 10854
rect 19272 10852 19296 10854
rect 19352 10852 19376 10854
rect 19432 10852 19456 10854
rect 19512 10852 19518 10854
rect 19210 10843 19518 10852
rect 26984 10908 27292 10917
rect 26984 10906 26990 10908
rect 27046 10906 27070 10908
rect 27126 10906 27150 10908
rect 27206 10906 27230 10908
rect 27286 10906 27292 10908
rect 27046 10854 27048 10906
rect 27228 10854 27230 10906
rect 26984 10852 26990 10854
rect 27046 10852 27070 10854
rect 27126 10852 27150 10854
rect 27206 10852 27230 10854
rect 27286 10852 27292 10854
rect 26984 10843 27292 10852
rect 19870 10364 20178 10373
rect 19870 10362 19876 10364
rect 19932 10362 19956 10364
rect 20012 10362 20036 10364
rect 20092 10362 20116 10364
rect 20172 10362 20178 10364
rect 19932 10310 19934 10362
rect 20114 10310 20116 10362
rect 19870 10308 19876 10310
rect 19932 10308 19956 10310
rect 20012 10308 20036 10310
rect 20092 10308 20116 10310
rect 20172 10308 20178 10310
rect 19870 10299 20178 10308
rect 27644 10364 27952 10373
rect 27644 10362 27650 10364
rect 27706 10362 27730 10364
rect 27786 10362 27810 10364
rect 27866 10362 27890 10364
rect 27946 10362 27952 10364
rect 27706 10310 27708 10362
rect 27888 10310 27890 10362
rect 27644 10308 27650 10310
rect 27706 10308 27730 10310
rect 27786 10308 27810 10310
rect 27866 10308 27890 10310
rect 27946 10308 27952 10310
rect 27644 10299 27952 10308
rect 19210 9820 19518 9829
rect 19210 9818 19216 9820
rect 19272 9818 19296 9820
rect 19352 9818 19376 9820
rect 19432 9818 19456 9820
rect 19512 9818 19518 9820
rect 19272 9766 19274 9818
rect 19454 9766 19456 9818
rect 19210 9764 19216 9766
rect 19272 9764 19296 9766
rect 19352 9764 19376 9766
rect 19432 9764 19456 9766
rect 19512 9764 19518 9766
rect 19210 9755 19518 9764
rect 26984 9820 27292 9829
rect 26984 9818 26990 9820
rect 27046 9818 27070 9820
rect 27126 9818 27150 9820
rect 27206 9818 27230 9820
rect 27286 9818 27292 9820
rect 27046 9766 27048 9818
rect 27228 9766 27230 9818
rect 26984 9764 26990 9766
rect 27046 9764 27070 9766
rect 27126 9764 27150 9766
rect 27206 9764 27230 9766
rect 27286 9764 27292 9766
rect 26984 9755 27292 9764
rect 19870 9276 20178 9285
rect 19870 9274 19876 9276
rect 19932 9274 19956 9276
rect 20012 9274 20036 9276
rect 20092 9274 20116 9276
rect 20172 9274 20178 9276
rect 19932 9222 19934 9274
rect 20114 9222 20116 9274
rect 19870 9220 19876 9222
rect 19932 9220 19956 9222
rect 20012 9220 20036 9222
rect 20092 9220 20116 9222
rect 20172 9220 20178 9222
rect 19870 9211 20178 9220
rect 27644 9276 27952 9285
rect 27644 9274 27650 9276
rect 27706 9274 27730 9276
rect 27786 9274 27810 9276
rect 27866 9274 27890 9276
rect 27946 9274 27952 9276
rect 27706 9222 27708 9274
rect 27888 9222 27890 9274
rect 27644 9220 27650 9222
rect 27706 9220 27730 9222
rect 27786 9220 27810 9222
rect 27866 9220 27890 9222
rect 27946 9220 27952 9222
rect 27644 9211 27952 9220
rect 19210 8732 19518 8741
rect 19210 8730 19216 8732
rect 19272 8730 19296 8732
rect 19352 8730 19376 8732
rect 19432 8730 19456 8732
rect 19512 8730 19518 8732
rect 19272 8678 19274 8730
rect 19454 8678 19456 8730
rect 19210 8676 19216 8678
rect 19272 8676 19296 8678
rect 19352 8676 19376 8678
rect 19432 8676 19456 8678
rect 19512 8676 19518 8678
rect 19210 8667 19518 8676
rect 26984 8732 27292 8741
rect 26984 8730 26990 8732
rect 27046 8730 27070 8732
rect 27126 8730 27150 8732
rect 27206 8730 27230 8732
rect 27286 8730 27292 8732
rect 27046 8678 27048 8730
rect 27228 8678 27230 8730
rect 26984 8676 26990 8678
rect 27046 8676 27070 8678
rect 27126 8676 27150 8678
rect 27206 8676 27230 8678
rect 27286 8676 27292 8678
rect 26984 8667 27292 8676
rect 19870 8188 20178 8197
rect 19870 8186 19876 8188
rect 19932 8186 19956 8188
rect 20012 8186 20036 8188
rect 20092 8186 20116 8188
rect 20172 8186 20178 8188
rect 19932 8134 19934 8186
rect 20114 8134 20116 8186
rect 19870 8132 19876 8134
rect 19932 8132 19956 8134
rect 20012 8132 20036 8134
rect 20092 8132 20116 8134
rect 20172 8132 20178 8134
rect 19870 8123 20178 8132
rect 27644 8188 27952 8197
rect 27644 8186 27650 8188
rect 27706 8186 27730 8188
rect 27786 8186 27810 8188
rect 27866 8186 27890 8188
rect 27946 8186 27952 8188
rect 27706 8134 27708 8186
rect 27888 8134 27890 8186
rect 27644 8132 27650 8134
rect 27706 8132 27730 8134
rect 27786 8132 27810 8134
rect 27866 8132 27890 8134
rect 27946 8132 27952 8134
rect 27644 8123 27952 8132
rect 19210 7644 19518 7653
rect 19210 7642 19216 7644
rect 19272 7642 19296 7644
rect 19352 7642 19376 7644
rect 19432 7642 19456 7644
rect 19512 7642 19518 7644
rect 19272 7590 19274 7642
rect 19454 7590 19456 7642
rect 19210 7588 19216 7590
rect 19272 7588 19296 7590
rect 19352 7588 19376 7590
rect 19432 7588 19456 7590
rect 19512 7588 19518 7590
rect 19210 7579 19518 7588
rect 26984 7644 27292 7653
rect 26984 7642 26990 7644
rect 27046 7642 27070 7644
rect 27126 7642 27150 7644
rect 27206 7642 27230 7644
rect 27286 7642 27292 7644
rect 27046 7590 27048 7642
rect 27228 7590 27230 7642
rect 26984 7588 26990 7590
rect 27046 7588 27070 7590
rect 27126 7588 27150 7590
rect 27206 7588 27230 7590
rect 27286 7588 27292 7590
rect 26984 7579 27292 7588
rect 19870 7100 20178 7109
rect 19870 7098 19876 7100
rect 19932 7098 19956 7100
rect 20012 7098 20036 7100
rect 20092 7098 20116 7100
rect 20172 7098 20178 7100
rect 19932 7046 19934 7098
rect 20114 7046 20116 7098
rect 19870 7044 19876 7046
rect 19932 7044 19956 7046
rect 20012 7044 20036 7046
rect 20092 7044 20116 7046
rect 20172 7044 20178 7046
rect 19870 7035 20178 7044
rect 27644 7100 27952 7109
rect 27644 7098 27650 7100
rect 27706 7098 27730 7100
rect 27786 7098 27810 7100
rect 27866 7098 27890 7100
rect 27946 7098 27952 7100
rect 27706 7046 27708 7098
rect 27888 7046 27890 7098
rect 27644 7044 27650 7046
rect 27706 7044 27730 7046
rect 27786 7044 27810 7046
rect 27866 7044 27890 7046
rect 27946 7044 27952 7046
rect 27644 7035 27952 7044
rect 17052 6886 17172 6914
rect 17052 1018 17080 6886
rect 19210 6556 19518 6565
rect 19210 6554 19216 6556
rect 19272 6554 19296 6556
rect 19352 6554 19376 6556
rect 19432 6554 19456 6556
rect 19512 6554 19518 6556
rect 19272 6502 19274 6554
rect 19454 6502 19456 6554
rect 19210 6500 19216 6502
rect 19272 6500 19296 6502
rect 19352 6500 19376 6502
rect 19432 6500 19456 6502
rect 19512 6500 19518 6502
rect 19210 6491 19518 6500
rect 26984 6556 27292 6565
rect 26984 6554 26990 6556
rect 27046 6554 27070 6556
rect 27126 6554 27150 6556
rect 27206 6554 27230 6556
rect 27286 6554 27292 6556
rect 27046 6502 27048 6554
rect 27228 6502 27230 6554
rect 26984 6500 26990 6502
rect 27046 6500 27070 6502
rect 27126 6500 27150 6502
rect 27206 6500 27230 6502
rect 27286 6500 27292 6502
rect 26984 6491 27292 6500
rect 19870 6012 20178 6021
rect 19870 6010 19876 6012
rect 19932 6010 19956 6012
rect 20012 6010 20036 6012
rect 20092 6010 20116 6012
rect 20172 6010 20178 6012
rect 19932 5958 19934 6010
rect 20114 5958 20116 6010
rect 19870 5956 19876 5958
rect 19932 5956 19956 5958
rect 20012 5956 20036 5958
rect 20092 5956 20116 5958
rect 20172 5956 20178 5958
rect 19870 5947 20178 5956
rect 27644 6012 27952 6021
rect 27644 6010 27650 6012
rect 27706 6010 27730 6012
rect 27786 6010 27810 6012
rect 27866 6010 27890 6012
rect 27946 6010 27952 6012
rect 27706 5958 27708 6010
rect 27888 5958 27890 6010
rect 27644 5956 27650 5958
rect 27706 5956 27730 5958
rect 27786 5956 27810 5958
rect 27866 5956 27890 5958
rect 27946 5956 27952 5958
rect 27644 5947 27952 5956
rect 19210 5468 19518 5477
rect 19210 5466 19216 5468
rect 19272 5466 19296 5468
rect 19352 5466 19376 5468
rect 19432 5466 19456 5468
rect 19512 5466 19518 5468
rect 19272 5414 19274 5466
rect 19454 5414 19456 5466
rect 19210 5412 19216 5414
rect 19272 5412 19296 5414
rect 19352 5412 19376 5414
rect 19432 5412 19456 5414
rect 19512 5412 19518 5414
rect 19210 5403 19518 5412
rect 26984 5468 27292 5477
rect 26984 5466 26990 5468
rect 27046 5466 27070 5468
rect 27126 5466 27150 5468
rect 27206 5466 27230 5468
rect 27286 5466 27292 5468
rect 27046 5414 27048 5466
rect 27228 5414 27230 5466
rect 26984 5412 26990 5414
rect 27046 5412 27070 5414
rect 27126 5412 27150 5414
rect 27206 5412 27230 5414
rect 27286 5412 27292 5414
rect 26984 5403 27292 5412
rect 19870 4924 20178 4933
rect 19870 4922 19876 4924
rect 19932 4922 19956 4924
rect 20012 4922 20036 4924
rect 20092 4922 20116 4924
rect 20172 4922 20178 4924
rect 19932 4870 19934 4922
rect 20114 4870 20116 4922
rect 19870 4868 19876 4870
rect 19932 4868 19956 4870
rect 20012 4868 20036 4870
rect 20092 4868 20116 4870
rect 20172 4868 20178 4870
rect 19870 4859 20178 4868
rect 27644 4924 27952 4933
rect 27644 4922 27650 4924
rect 27706 4922 27730 4924
rect 27786 4922 27810 4924
rect 27866 4922 27890 4924
rect 27946 4922 27952 4924
rect 27706 4870 27708 4922
rect 27888 4870 27890 4922
rect 27644 4868 27650 4870
rect 27706 4868 27730 4870
rect 27786 4868 27810 4870
rect 27866 4868 27890 4870
rect 27946 4868 27952 4870
rect 27644 4859 27952 4868
rect 19210 4380 19518 4389
rect 19210 4378 19216 4380
rect 19272 4378 19296 4380
rect 19352 4378 19376 4380
rect 19432 4378 19456 4380
rect 19512 4378 19518 4380
rect 19272 4326 19274 4378
rect 19454 4326 19456 4378
rect 19210 4324 19216 4326
rect 19272 4324 19296 4326
rect 19352 4324 19376 4326
rect 19432 4324 19456 4326
rect 19512 4324 19518 4326
rect 19210 4315 19518 4324
rect 26984 4380 27292 4389
rect 26984 4378 26990 4380
rect 27046 4378 27070 4380
rect 27126 4378 27150 4380
rect 27206 4378 27230 4380
rect 27286 4378 27292 4380
rect 27046 4326 27048 4378
rect 27228 4326 27230 4378
rect 26984 4324 26990 4326
rect 27046 4324 27070 4326
rect 27126 4324 27150 4326
rect 27206 4324 27230 4326
rect 27286 4324 27292 4326
rect 26984 4315 27292 4324
rect 19870 3836 20178 3845
rect 19870 3834 19876 3836
rect 19932 3834 19956 3836
rect 20012 3834 20036 3836
rect 20092 3834 20116 3836
rect 20172 3834 20178 3836
rect 19932 3782 19934 3834
rect 20114 3782 20116 3834
rect 19870 3780 19876 3782
rect 19932 3780 19956 3782
rect 20012 3780 20036 3782
rect 20092 3780 20116 3782
rect 20172 3780 20178 3782
rect 19870 3771 20178 3780
rect 27644 3836 27952 3845
rect 27644 3834 27650 3836
rect 27706 3834 27730 3836
rect 27786 3834 27810 3836
rect 27866 3834 27890 3836
rect 27946 3834 27952 3836
rect 27706 3782 27708 3834
rect 27888 3782 27890 3834
rect 27644 3780 27650 3782
rect 27706 3780 27730 3782
rect 27786 3780 27810 3782
rect 27866 3780 27890 3782
rect 27946 3780 27952 3782
rect 27644 3771 27952 3780
rect 19210 3292 19518 3301
rect 19210 3290 19216 3292
rect 19272 3290 19296 3292
rect 19352 3290 19376 3292
rect 19432 3290 19456 3292
rect 19512 3290 19518 3292
rect 19272 3238 19274 3290
rect 19454 3238 19456 3290
rect 19210 3236 19216 3238
rect 19272 3236 19296 3238
rect 19352 3236 19376 3238
rect 19432 3236 19456 3238
rect 19512 3236 19518 3238
rect 19210 3227 19518 3236
rect 26984 3292 27292 3301
rect 26984 3290 26990 3292
rect 27046 3290 27070 3292
rect 27126 3290 27150 3292
rect 27206 3290 27230 3292
rect 27286 3290 27292 3292
rect 27046 3238 27048 3290
rect 27228 3238 27230 3290
rect 26984 3236 26990 3238
rect 27046 3236 27070 3238
rect 27126 3236 27150 3238
rect 27206 3236 27230 3238
rect 27286 3236 27292 3238
rect 26984 3227 27292 3236
rect 19870 2748 20178 2757
rect 19870 2746 19876 2748
rect 19932 2746 19956 2748
rect 20012 2746 20036 2748
rect 20092 2746 20116 2748
rect 20172 2746 20178 2748
rect 19932 2694 19934 2746
rect 20114 2694 20116 2746
rect 19870 2692 19876 2694
rect 19932 2692 19956 2694
rect 20012 2692 20036 2694
rect 20092 2692 20116 2694
rect 20172 2692 20178 2694
rect 19870 2683 20178 2692
rect 27644 2748 27952 2757
rect 27644 2746 27650 2748
rect 27706 2746 27730 2748
rect 27786 2746 27810 2748
rect 27866 2746 27890 2748
rect 27946 2746 27952 2748
rect 27706 2694 27708 2746
rect 27888 2694 27890 2746
rect 27644 2692 27650 2694
rect 27706 2692 27730 2694
rect 27786 2692 27810 2694
rect 27866 2692 27890 2694
rect 27946 2692 27952 2694
rect 27644 2683 27952 2692
rect 19210 2204 19518 2213
rect 19210 2202 19216 2204
rect 19272 2202 19296 2204
rect 19352 2202 19376 2204
rect 19432 2202 19456 2204
rect 19512 2202 19518 2204
rect 19272 2150 19274 2202
rect 19454 2150 19456 2202
rect 19210 2148 19216 2150
rect 19272 2148 19296 2150
rect 19352 2148 19376 2150
rect 19432 2148 19456 2150
rect 19512 2148 19518 2150
rect 19210 2139 19518 2148
rect 26984 2204 27292 2213
rect 26984 2202 26990 2204
rect 27046 2202 27070 2204
rect 27126 2202 27150 2204
rect 27206 2202 27230 2204
rect 27286 2202 27292 2204
rect 27046 2150 27048 2202
rect 27228 2150 27230 2202
rect 26984 2148 26990 2150
rect 27046 2148 27070 2150
rect 27126 2148 27150 2150
rect 27206 2148 27230 2150
rect 27286 2148 27292 2150
rect 26984 2139 27292 2148
rect 19870 1660 20178 1669
rect 19870 1658 19876 1660
rect 19932 1658 19956 1660
rect 20012 1658 20036 1660
rect 20092 1658 20116 1660
rect 20172 1658 20178 1660
rect 19932 1606 19934 1658
rect 20114 1606 20116 1658
rect 19870 1604 19876 1606
rect 19932 1604 19956 1606
rect 20012 1604 20036 1606
rect 20092 1604 20116 1606
rect 20172 1604 20178 1606
rect 19870 1595 20178 1604
rect 27644 1660 27952 1669
rect 27644 1658 27650 1660
rect 27706 1658 27730 1660
rect 27786 1658 27810 1660
rect 27866 1658 27890 1660
rect 27946 1658 27952 1660
rect 27706 1606 27708 1658
rect 27888 1606 27890 1658
rect 27644 1604 27650 1606
rect 27706 1604 27730 1606
rect 27786 1604 27810 1606
rect 27866 1604 27890 1606
rect 27946 1604 27952 1606
rect 27644 1595 27952 1604
rect 19210 1116 19518 1125
rect 19210 1114 19216 1116
rect 19272 1114 19296 1116
rect 19352 1114 19376 1116
rect 19432 1114 19456 1116
rect 19512 1114 19518 1116
rect 19272 1062 19274 1114
rect 19454 1062 19456 1114
rect 19210 1060 19216 1062
rect 19272 1060 19296 1062
rect 19352 1060 19376 1062
rect 19432 1060 19456 1062
rect 19512 1060 19518 1062
rect 19210 1051 19518 1060
rect 26984 1116 27292 1125
rect 26984 1114 26990 1116
rect 27046 1114 27070 1116
rect 27126 1114 27150 1116
rect 27206 1114 27230 1116
rect 27286 1114 27292 1116
rect 27046 1062 27048 1114
rect 27228 1062 27230 1114
rect 26984 1060 26990 1062
rect 27046 1060 27070 1062
rect 27126 1060 27150 1062
rect 27206 1060 27230 1062
rect 27286 1060 27292 1062
rect 26984 1051 27292 1060
rect 17040 1012 17092 1018
rect 17040 954 17092 960
rect 16120 944 16172 950
rect 16120 886 16172 892
rect 16764 944 16816 950
rect 16764 886 16816 892
rect 7104 808 7156 814
rect 7104 750 7156 756
rect 9036 808 9088 814
rect 9036 750 9088 756
rect 11612 808 11664 814
rect 11612 750 11664 756
rect 12440 808 12492 814
rect 12440 750 12492 756
rect 12900 808 12952 814
rect 12900 750 12952 756
rect 13544 808 13596 814
rect 13544 750 13596 756
rect 14188 808 14240 814
rect 14188 750 14240 756
rect 14832 808 14884 814
rect 14832 750 14884 756
rect 15476 808 15528 814
rect 15476 750 15528 756
rect 4322 572 4630 581
rect 4322 570 4328 572
rect 4384 570 4408 572
rect 4464 570 4488 572
rect 4544 570 4568 572
rect 4624 570 4630 572
rect 4384 518 4386 570
rect 4566 518 4568 570
rect 4322 516 4328 518
rect 4384 516 4408 518
rect 4464 516 4488 518
rect 4544 516 4568 518
rect 4624 516 4630 518
rect 4322 507 4630 516
rect 7116 400 7144 750
rect 9048 400 9076 750
rect 11624 400 11652 750
rect 12096 572 12404 581
rect 12096 570 12102 572
rect 12158 570 12182 572
rect 12238 570 12262 572
rect 12318 570 12342 572
rect 12398 570 12404 572
rect 12158 518 12160 570
rect 12340 518 12342 570
rect 12096 516 12102 518
rect 12158 516 12182 518
rect 12238 516 12262 518
rect 12318 516 12342 518
rect 12398 516 12404 518
rect 12096 507 12404 516
rect 12452 474 12480 750
rect 12164 468 12216 474
rect 12440 468 12492 474
rect 12216 428 12296 456
rect 12164 410 12216 416
rect 12268 400 12296 428
rect 12440 410 12492 416
rect 12912 400 12940 750
rect 13556 400 13584 750
rect 14200 400 14228 750
rect 14844 400 14872 750
rect 15488 400 15516 750
rect 16132 400 16160 886
rect 16764 808 16816 814
rect 16764 750 16816 756
rect 17408 808 17460 814
rect 17408 750 17460 756
rect 18052 808 18104 814
rect 18052 750 18104 756
rect 18696 808 18748 814
rect 18696 750 18748 756
rect 19800 808 19852 814
rect 19800 750 19852 756
rect 16776 400 16804 750
rect 17420 400 17448 750
rect 18064 400 18092 750
rect 18708 400 18736 750
rect 19812 456 19840 750
rect 19870 572 20178 581
rect 19870 570 19876 572
rect 19932 570 19956 572
rect 20012 570 20036 572
rect 20092 570 20116 572
rect 20172 570 20178 572
rect 19932 518 19934 570
rect 20114 518 20116 570
rect 19870 516 19876 518
rect 19932 516 19956 518
rect 20012 516 20036 518
rect 20092 516 20116 518
rect 20172 516 20178 518
rect 19870 507 20178 516
rect 27644 572 27952 581
rect 27644 570 27650 572
rect 27706 570 27730 572
rect 27786 570 27810 572
rect 27866 570 27890 572
rect 27946 570 27952 572
rect 27706 518 27708 570
rect 27888 518 27890 570
rect 27644 516 27650 518
rect 27706 516 27730 518
rect 27786 516 27810 518
rect 27866 516 27890 518
rect 27946 516 27952 518
rect 27644 507 27952 516
rect 19812 428 20024 456
rect 19996 400 20024 428
rect 18 0 74 400
rect 662 0 718 400
rect 1306 0 1362 400
rect 1950 0 2006 400
rect 2594 0 2650 400
rect 3238 0 3294 400
rect 3882 0 3938 400
rect 4526 0 4582 400
rect 5170 0 5226 400
rect 5814 0 5870 400
rect 6458 0 6514 400
rect 7102 0 7158 400
rect 7746 0 7802 400
rect 8390 0 8446 400
rect 9034 0 9090 400
rect 9678 0 9734 400
rect 10322 0 10378 400
rect 10966 0 11022 400
rect 11610 0 11666 400
rect 12254 0 12310 400
rect 12898 0 12954 400
rect 13542 0 13598 400
rect 14186 0 14242 400
rect 14830 0 14886 400
rect 15474 0 15530 400
rect 16118 0 16174 400
rect 16762 0 16818 400
rect 17406 0 17462 400
rect 18050 0 18106 400
rect 18694 0 18750 400
rect 19982 0 20038 400
<< via2 >>
rect 4328 19066 4384 19068
rect 4408 19066 4464 19068
rect 4488 19066 4544 19068
rect 4568 19066 4624 19068
rect 4328 19014 4374 19066
rect 4374 19014 4384 19066
rect 4408 19014 4438 19066
rect 4438 19014 4450 19066
rect 4450 19014 4464 19066
rect 4488 19014 4502 19066
rect 4502 19014 4514 19066
rect 4514 19014 4544 19066
rect 4568 19014 4578 19066
rect 4578 19014 4624 19066
rect 4328 19012 4384 19014
rect 4408 19012 4464 19014
rect 4488 19012 4544 19014
rect 4568 19012 4624 19014
rect 12102 19066 12158 19068
rect 12182 19066 12238 19068
rect 12262 19066 12318 19068
rect 12342 19066 12398 19068
rect 12102 19014 12148 19066
rect 12148 19014 12158 19066
rect 12182 19014 12212 19066
rect 12212 19014 12224 19066
rect 12224 19014 12238 19066
rect 12262 19014 12276 19066
rect 12276 19014 12288 19066
rect 12288 19014 12318 19066
rect 12342 19014 12352 19066
rect 12352 19014 12398 19066
rect 12102 19012 12158 19014
rect 12182 19012 12238 19014
rect 12262 19012 12318 19014
rect 12342 19012 12398 19014
rect 3668 18522 3724 18524
rect 3748 18522 3804 18524
rect 3828 18522 3884 18524
rect 3908 18522 3964 18524
rect 3668 18470 3714 18522
rect 3714 18470 3724 18522
rect 3748 18470 3778 18522
rect 3778 18470 3790 18522
rect 3790 18470 3804 18522
rect 3828 18470 3842 18522
rect 3842 18470 3854 18522
rect 3854 18470 3884 18522
rect 3908 18470 3918 18522
rect 3918 18470 3964 18522
rect 3668 18468 3724 18470
rect 3748 18468 3804 18470
rect 3828 18468 3884 18470
rect 3908 18468 3964 18470
rect 11442 18522 11498 18524
rect 11522 18522 11578 18524
rect 11602 18522 11658 18524
rect 11682 18522 11738 18524
rect 11442 18470 11488 18522
rect 11488 18470 11498 18522
rect 11522 18470 11552 18522
rect 11552 18470 11564 18522
rect 11564 18470 11578 18522
rect 11602 18470 11616 18522
rect 11616 18470 11628 18522
rect 11628 18470 11658 18522
rect 11682 18470 11692 18522
rect 11692 18470 11738 18522
rect 11442 18468 11498 18470
rect 11522 18468 11578 18470
rect 11602 18468 11658 18470
rect 11682 18468 11738 18470
rect 846 18400 902 18456
rect 4328 17978 4384 17980
rect 4408 17978 4464 17980
rect 4488 17978 4544 17980
rect 4568 17978 4624 17980
rect 4328 17926 4374 17978
rect 4374 17926 4384 17978
rect 4408 17926 4438 17978
rect 4438 17926 4450 17978
rect 4450 17926 4464 17978
rect 4488 17926 4502 17978
rect 4502 17926 4514 17978
rect 4514 17926 4544 17978
rect 4568 17926 4578 17978
rect 4578 17926 4624 17978
rect 4328 17924 4384 17926
rect 4408 17924 4464 17926
rect 4488 17924 4544 17926
rect 4568 17924 4624 17926
rect 12102 17978 12158 17980
rect 12182 17978 12238 17980
rect 12262 17978 12318 17980
rect 12342 17978 12398 17980
rect 12102 17926 12148 17978
rect 12148 17926 12158 17978
rect 12182 17926 12212 17978
rect 12212 17926 12224 17978
rect 12224 17926 12238 17978
rect 12262 17926 12276 17978
rect 12276 17926 12288 17978
rect 12288 17926 12318 17978
rect 12342 17926 12352 17978
rect 12352 17926 12398 17978
rect 12102 17924 12158 17926
rect 12182 17924 12238 17926
rect 12262 17924 12318 17926
rect 12342 17924 12398 17926
rect 3668 17434 3724 17436
rect 3748 17434 3804 17436
rect 3828 17434 3884 17436
rect 3908 17434 3964 17436
rect 3668 17382 3714 17434
rect 3714 17382 3724 17434
rect 3748 17382 3778 17434
rect 3778 17382 3790 17434
rect 3790 17382 3804 17434
rect 3828 17382 3842 17434
rect 3842 17382 3854 17434
rect 3854 17382 3884 17434
rect 3908 17382 3918 17434
rect 3918 17382 3964 17434
rect 3668 17380 3724 17382
rect 3748 17380 3804 17382
rect 3828 17380 3884 17382
rect 3908 17380 3964 17382
rect 11442 17434 11498 17436
rect 11522 17434 11578 17436
rect 11602 17434 11658 17436
rect 11682 17434 11738 17436
rect 11442 17382 11488 17434
rect 11488 17382 11498 17434
rect 11522 17382 11552 17434
rect 11552 17382 11564 17434
rect 11564 17382 11578 17434
rect 11602 17382 11616 17434
rect 11616 17382 11628 17434
rect 11628 17382 11658 17434
rect 11682 17382 11692 17434
rect 11692 17382 11738 17434
rect 11442 17380 11498 17382
rect 11522 17380 11578 17382
rect 11602 17380 11658 17382
rect 11682 17380 11738 17382
rect 4328 16890 4384 16892
rect 4408 16890 4464 16892
rect 4488 16890 4544 16892
rect 4568 16890 4624 16892
rect 4328 16838 4374 16890
rect 4374 16838 4384 16890
rect 4408 16838 4438 16890
rect 4438 16838 4450 16890
rect 4450 16838 4464 16890
rect 4488 16838 4502 16890
rect 4502 16838 4514 16890
rect 4514 16838 4544 16890
rect 4568 16838 4578 16890
rect 4578 16838 4624 16890
rect 4328 16836 4384 16838
rect 4408 16836 4464 16838
rect 4488 16836 4544 16838
rect 4568 16836 4624 16838
rect 12102 16890 12158 16892
rect 12182 16890 12238 16892
rect 12262 16890 12318 16892
rect 12342 16890 12398 16892
rect 12102 16838 12148 16890
rect 12148 16838 12158 16890
rect 12182 16838 12212 16890
rect 12212 16838 12224 16890
rect 12224 16838 12238 16890
rect 12262 16838 12276 16890
rect 12276 16838 12288 16890
rect 12288 16838 12318 16890
rect 12342 16838 12352 16890
rect 12352 16838 12398 16890
rect 12102 16836 12158 16838
rect 12182 16836 12238 16838
rect 12262 16836 12318 16838
rect 12342 16836 12398 16838
rect 14370 17720 14426 17776
rect 3668 16346 3724 16348
rect 3748 16346 3804 16348
rect 3828 16346 3884 16348
rect 3908 16346 3964 16348
rect 3668 16294 3714 16346
rect 3714 16294 3724 16346
rect 3748 16294 3778 16346
rect 3778 16294 3790 16346
rect 3790 16294 3804 16346
rect 3828 16294 3842 16346
rect 3842 16294 3854 16346
rect 3854 16294 3884 16346
rect 3908 16294 3918 16346
rect 3918 16294 3964 16346
rect 3668 16292 3724 16294
rect 3748 16292 3804 16294
rect 3828 16292 3884 16294
rect 3908 16292 3964 16294
rect 11442 16346 11498 16348
rect 11522 16346 11578 16348
rect 11602 16346 11658 16348
rect 11682 16346 11738 16348
rect 11442 16294 11488 16346
rect 11488 16294 11498 16346
rect 11522 16294 11552 16346
rect 11552 16294 11564 16346
rect 11564 16294 11578 16346
rect 11602 16294 11616 16346
rect 11616 16294 11628 16346
rect 11628 16294 11658 16346
rect 11682 16294 11692 16346
rect 11692 16294 11738 16346
rect 11442 16292 11498 16294
rect 11522 16292 11578 16294
rect 11602 16292 11658 16294
rect 11682 16292 11738 16294
rect 4328 15802 4384 15804
rect 4408 15802 4464 15804
rect 4488 15802 4544 15804
rect 4568 15802 4624 15804
rect 4328 15750 4374 15802
rect 4374 15750 4384 15802
rect 4408 15750 4438 15802
rect 4438 15750 4450 15802
rect 4450 15750 4464 15802
rect 4488 15750 4502 15802
rect 4502 15750 4514 15802
rect 4514 15750 4544 15802
rect 4568 15750 4578 15802
rect 4578 15750 4624 15802
rect 4328 15748 4384 15750
rect 4408 15748 4464 15750
rect 4488 15748 4544 15750
rect 4568 15748 4624 15750
rect 12102 15802 12158 15804
rect 12182 15802 12238 15804
rect 12262 15802 12318 15804
rect 12342 15802 12398 15804
rect 12102 15750 12148 15802
rect 12148 15750 12158 15802
rect 12182 15750 12212 15802
rect 12212 15750 12224 15802
rect 12224 15750 12238 15802
rect 12262 15750 12276 15802
rect 12276 15750 12288 15802
rect 12288 15750 12318 15802
rect 12342 15750 12352 15802
rect 12352 15750 12398 15802
rect 12102 15748 12158 15750
rect 12182 15748 12238 15750
rect 12262 15748 12318 15750
rect 12342 15748 12398 15750
rect 3668 15258 3724 15260
rect 3748 15258 3804 15260
rect 3828 15258 3884 15260
rect 3908 15258 3964 15260
rect 3668 15206 3714 15258
rect 3714 15206 3724 15258
rect 3748 15206 3778 15258
rect 3778 15206 3790 15258
rect 3790 15206 3804 15258
rect 3828 15206 3842 15258
rect 3842 15206 3854 15258
rect 3854 15206 3884 15258
rect 3908 15206 3918 15258
rect 3918 15206 3964 15258
rect 3668 15204 3724 15206
rect 3748 15204 3804 15206
rect 3828 15204 3884 15206
rect 3908 15204 3964 15206
rect 11442 15258 11498 15260
rect 11522 15258 11578 15260
rect 11602 15258 11658 15260
rect 11682 15258 11738 15260
rect 11442 15206 11488 15258
rect 11488 15206 11498 15258
rect 11522 15206 11552 15258
rect 11552 15206 11564 15258
rect 11564 15206 11578 15258
rect 11602 15206 11616 15258
rect 11616 15206 11628 15258
rect 11628 15206 11658 15258
rect 11682 15206 11692 15258
rect 11692 15206 11738 15258
rect 11442 15204 11498 15206
rect 11522 15204 11578 15206
rect 11602 15204 11658 15206
rect 11682 15204 11738 15206
rect 4328 14714 4384 14716
rect 4408 14714 4464 14716
rect 4488 14714 4544 14716
rect 4568 14714 4624 14716
rect 4328 14662 4374 14714
rect 4374 14662 4384 14714
rect 4408 14662 4438 14714
rect 4438 14662 4450 14714
rect 4450 14662 4464 14714
rect 4488 14662 4502 14714
rect 4502 14662 4514 14714
rect 4514 14662 4544 14714
rect 4568 14662 4578 14714
rect 4578 14662 4624 14714
rect 4328 14660 4384 14662
rect 4408 14660 4464 14662
rect 4488 14660 4544 14662
rect 4568 14660 4624 14662
rect 12102 14714 12158 14716
rect 12182 14714 12238 14716
rect 12262 14714 12318 14716
rect 12342 14714 12398 14716
rect 12102 14662 12148 14714
rect 12148 14662 12158 14714
rect 12182 14662 12212 14714
rect 12212 14662 12224 14714
rect 12224 14662 12238 14714
rect 12262 14662 12276 14714
rect 12276 14662 12288 14714
rect 12288 14662 12318 14714
rect 12342 14662 12352 14714
rect 12352 14662 12398 14714
rect 12102 14660 12158 14662
rect 12182 14660 12238 14662
rect 12262 14660 12318 14662
rect 12342 14660 12398 14662
rect 15014 17740 15070 17776
rect 15014 17720 15016 17740
rect 15016 17720 15068 17740
rect 15068 17720 15070 17740
rect 19876 19066 19932 19068
rect 19956 19066 20012 19068
rect 20036 19066 20092 19068
rect 20116 19066 20172 19068
rect 19876 19014 19922 19066
rect 19922 19014 19932 19066
rect 19956 19014 19986 19066
rect 19986 19014 19998 19066
rect 19998 19014 20012 19066
rect 20036 19014 20050 19066
rect 20050 19014 20062 19066
rect 20062 19014 20092 19066
rect 20116 19014 20126 19066
rect 20126 19014 20172 19066
rect 19876 19012 19932 19014
rect 19956 19012 20012 19014
rect 20036 19012 20092 19014
rect 20116 19012 20172 19014
rect 27650 19066 27706 19068
rect 27730 19066 27786 19068
rect 27810 19066 27866 19068
rect 27890 19066 27946 19068
rect 27650 19014 27696 19066
rect 27696 19014 27706 19066
rect 27730 19014 27760 19066
rect 27760 19014 27772 19066
rect 27772 19014 27786 19066
rect 27810 19014 27824 19066
rect 27824 19014 27836 19066
rect 27836 19014 27866 19066
rect 27890 19014 27900 19066
rect 27900 19014 27946 19066
rect 27650 19012 27706 19014
rect 27730 19012 27786 19014
rect 27810 19012 27866 19014
rect 27890 19012 27946 19014
rect 3668 14170 3724 14172
rect 3748 14170 3804 14172
rect 3828 14170 3884 14172
rect 3908 14170 3964 14172
rect 3668 14118 3714 14170
rect 3714 14118 3724 14170
rect 3748 14118 3778 14170
rect 3778 14118 3790 14170
rect 3790 14118 3804 14170
rect 3828 14118 3842 14170
rect 3842 14118 3854 14170
rect 3854 14118 3884 14170
rect 3908 14118 3918 14170
rect 3918 14118 3964 14170
rect 3668 14116 3724 14118
rect 3748 14116 3804 14118
rect 3828 14116 3884 14118
rect 3908 14116 3964 14118
rect 11442 14170 11498 14172
rect 11522 14170 11578 14172
rect 11602 14170 11658 14172
rect 11682 14170 11738 14172
rect 11442 14118 11488 14170
rect 11488 14118 11498 14170
rect 11522 14118 11552 14170
rect 11552 14118 11564 14170
rect 11564 14118 11578 14170
rect 11602 14118 11616 14170
rect 11616 14118 11628 14170
rect 11628 14118 11658 14170
rect 11682 14118 11692 14170
rect 11692 14118 11738 14170
rect 11442 14116 11498 14118
rect 11522 14116 11578 14118
rect 11602 14116 11658 14118
rect 11682 14116 11738 14118
rect 19216 18522 19272 18524
rect 19296 18522 19352 18524
rect 19376 18522 19432 18524
rect 19456 18522 19512 18524
rect 19216 18470 19262 18522
rect 19262 18470 19272 18522
rect 19296 18470 19326 18522
rect 19326 18470 19338 18522
rect 19338 18470 19352 18522
rect 19376 18470 19390 18522
rect 19390 18470 19402 18522
rect 19402 18470 19432 18522
rect 19456 18470 19466 18522
rect 19466 18470 19512 18522
rect 19216 18468 19272 18470
rect 19296 18468 19352 18470
rect 19376 18468 19432 18470
rect 19456 18468 19512 18470
rect 26990 18522 27046 18524
rect 27070 18522 27126 18524
rect 27150 18522 27206 18524
rect 27230 18522 27286 18524
rect 26990 18470 27036 18522
rect 27036 18470 27046 18522
rect 27070 18470 27100 18522
rect 27100 18470 27112 18522
rect 27112 18470 27126 18522
rect 27150 18470 27164 18522
rect 27164 18470 27176 18522
rect 27176 18470 27206 18522
rect 27230 18470 27240 18522
rect 27240 18470 27286 18522
rect 26990 18468 27046 18470
rect 27070 18468 27126 18470
rect 27150 18468 27206 18470
rect 27230 18468 27286 18470
rect 19876 17978 19932 17980
rect 19956 17978 20012 17980
rect 20036 17978 20092 17980
rect 20116 17978 20172 17980
rect 19876 17926 19922 17978
rect 19922 17926 19932 17978
rect 19956 17926 19986 17978
rect 19986 17926 19998 17978
rect 19998 17926 20012 17978
rect 20036 17926 20050 17978
rect 20050 17926 20062 17978
rect 20062 17926 20092 17978
rect 20116 17926 20126 17978
rect 20126 17926 20172 17978
rect 19876 17924 19932 17926
rect 19956 17924 20012 17926
rect 20036 17924 20092 17926
rect 20116 17924 20172 17926
rect 27650 17978 27706 17980
rect 27730 17978 27786 17980
rect 27810 17978 27866 17980
rect 27890 17978 27946 17980
rect 27650 17926 27696 17978
rect 27696 17926 27706 17978
rect 27730 17926 27760 17978
rect 27760 17926 27772 17978
rect 27772 17926 27786 17978
rect 27810 17926 27824 17978
rect 27824 17926 27836 17978
rect 27836 17926 27866 17978
rect 27890 17926 27900 17978
rect 27900 17926 27946 17978
rect 27650 17924 27706 17926
rect 27730 17924 27786 17926
rect 27810 17924 27866 17926
rect 27890 17924 27946 17926
rect 4328 13626 4384 13628
rect 4408 13626 4464 13628
rect 4488 13626 4544 13628
rect 4568 13626 4624 13628
rect 4328 13574 4374 13626
rect 4374 13574 4384 13626
rect 4408 13574 4438 13626
rect 4438 13574 4450 13626
rect 4450 13574 4464 13626
rect 4488 13574 4502 13626
rect 4502 13574 4514 13626
rect 4514 13574 4544 13626
rect 4568 13574 4578 13626
rect 4578 13574 4624 13626
rect 4328 13572 4384 13574
rect 4408 13572 4464 13574
rect 4488 13572 4544 13574
rect 4568 13572 4624 13574
rect 12102 13626 12158 13628
rect 12182 13626 12238 13628
rect 12262 13626 12318 13628
rect 12342 13626 12398 13628
rect 12102 13574 12148 13626
rect 12148 13574 12158 13626
rect 12182 13574 12212 13626
rect 12212 13574 12224 13626
rect 12224 13574 12238 13626
rect 12262 13574 12276 13626
rect 12276 13574 12288 13626
rect 12288 13574 12318 13626
rect 12342 13574 12352 13626
rect 12352 13574 12398 13626
rect 12102 13572 12158 13574
rect 12182 13572 12238 13574
rect 12262 13572 12318 13574
rect 12342 13572 12398 13574
rect 3668 13082 3724 13084
rect 3748 13082 3804 13084
rect 3828 13082 3884 13084
rect 3908 13082 3964 13084
rect 3668 13030 3714 13082
rect 3714 13030 3724 13082
rect 3748 13030 3778 13082
rect 3778 13030 3790 13082
rect 3790 13030 3804 13082
rect 3828 13030 3842 13082
rect 3842 13030 3854 13082
rect 3854 13030 3884 13082
rect 3908 13030 3918 13082
rect 3918 13030 3964 13082
rect 3668 13028 3724 13030
rect 3748 13028 3804 13030
rect 3828 13028 3884 13030
rect 3908 13028 3964 13030
rect 11442 13082 11498 13084
rect 11522 13082 11578 13084
rect 11602 13082 11658 13084
rect 11682 13082 11738 13084
rect 11442 13030 11488 13082
rect 11488 13030 11498 13082
rect 11522 13030 11552 13082
rect 11552 13030 11564 13082
rect 11564 13030 11578 13082
rect 11602 13030 11616 13082
rect 11616 13030 11628 13082
rect 11628 13030 11658 13082
rect 11682 13030 11692 13082
rect 11692 13030 11738 13082
rect 11442 13028 11498 13030
rect 11522 13028 11578 13030
rect 11602 13028 11658 13030
rect 11682 13028 11738 13030
rect 4328 12538 4384 12540
rect 4408 12538 4464 12540
rect 4488 12538 4544 12540
rect 4568 12538 4624 12540
rect 4328 12486 4374 12538
rect 4374 12486 4384 12538
rect 4408 12486 4438 12538
rect 4438 12486 4450 12538
rect 4450 12486 4464 12538
rect 4488 12486 4502 12538
rect 4502 12486 4514 12538
rect 4514 12486 4544 12538
rect 4568 12486 4578 12538
rect 4578 12486 4624 12538
rect 4328 12484 4384 12486
rect 4408 12484 4464 12486
rect 4488 12484 4544 12486
rect 4568 12484 4624 12486
rect 12102 12538 12158 12540
rect 12182 12538 12238 12540
rect 12262 12538 12318 12540
rect 12342 12538 12398 12540
rect 12102 12486 12148 12538
rect 12148 12486 12158 12538
rect 12182 12486 12212 12538
rect 12212 12486 12224 12538
rect 12224 12486 12238 12538
rect 12262 12486 12276 12538
rect 12276 12486 12288 12538
rect 12288 12486 12318 12538
rect 12342 12486 12352 12538
rect 12352 12486 12398 12538
rect 12102 12484 12158 12486
rect 12182 12484 12238 12486
rect 12262 12484 12318 12486
rect 12342 12484 12398 12486
rect 3668 11994 3724 11996
rect 3748 11994 3804 11996
rect 3828 11994 3884 11996
rect 3908 11994 3964 11996
rect 3668 11942 3714 11994
rect 3714 11942 3724 11994
rect 3748 11942 3778 11994
rect 3778 11942 3790 11994
rect 3790 11942 3804 11994
rect 3828 11942 3842 11994
rect 3842 11942 3854 11994
rect 3854 11942 3884 11994
rect 3908 11942 3918 11994
rect 3918 11942 3964 11994
rect 3668 11940 3724 11942
rect 3748 11940 3804 11942
rect 3828 11940 3884 11942
rect 3908 11940 3964 11942
rect 11442 11994 11498 11996
rect 11522 11994 11578 11996
rect 11602 11994 11658 11996
rect 11682 11994 11738 11996
rect 11442 11942 11488 11994
rect 11488 11942 11498 11994
rect 11522 11942 11552 11994
rect 11552 11942 11564 11994
rect 11564 11942 11578 11994
rect 11602 11942 11616 11994
rect 11616 11942 11628 11994
rect 11628 11942 11658 11994
rect 11682 11942 11692 11994
rect 11692 11942 11738 11994
rect 11442 11940 11498 11942
rect 11522 11940 11578 11942
rect 11602 11940 11658 11942
rect 11682 11940 11738 11942
rect 4328 11450 4384 11452
rect 4408 11450 4464 11452
rect 4488 11450 4544 11452
rect 4568 11450 4624 11452
rect 4328 11398 4374 11450
rect 4374 11398 4384 11450
rect 4408 11398 4438 11450
rect 4438 11398 4450 11450
rect 4450 11398 4464 11450
rect 4488 11398 4502 11450
rect 4502 11398 4514 11450
rect 4514 11398 4544 11450
rect 4568 11398 4578 11450
rect 4578 11398 4624 11450
rect 4328 11396 4384 11398
rect 4408 11396 4464 11398
rect 4488 11396 4544 11398
rect 4568 11396 4624 11398
rect 12102 11450 12158 11452
rect 12182 11450 12238 11452
rect 12262 11450 12318 11452
rect 12342 11450 12398 11452
rect 12102 11398 12148 11450
rect 12148 11398 12158 11450
rect 12182 11398 12212 11450
rect 12212 11398 12224 11450
rect 12224 11398 12238 11450
rect 12262 11398 12276 11450
rect 12276 11398 12288 11450
rect 12288 11398 12318 11450
rect 12342 11398 12352 11450
rect 12352 11398 12398 11450
rect 12102 11396 12158 11398
rect 12182 11396 12238 11398
rect 12262 11396 12318 11398
rect 12342 11396 12398 11398
rect 3668 10906 3724 10908
rect 3748 10906 3804 10908
rect 3828 10906 3884 10908
rect 3908 10906 3964 10908
rect 3668 10854 3714 10906
rect 3714 10854 3724 10906
rect 3748 10854 3778 10906
rect 3778 10854 3790 10906
rect 3790 10854 3804 10906
rect 3828 10854 3842 10906
rect 3842 10854 3854 10906
rect 3854 10854 3884 10906
rect 3908 10854 3918 10906
rect 3918 10854 3964 10906
rect 3668 10852 3724 10854
rect 3748 10852 3804 10854
rect 3828 10852 3884 10854
rect 3908 10852 3964 10854
rect 11442 10906 11498 10908
rect 11522 10906 11578 10908
rect 11602 10906 11658 10908
rect 11682 10906 11738 10908
rect 11442 10854 11488 10906
rect 11488 10854 11498 10906
rect 11522 10854 11552 10906
rect 11552 10854 11564 10906
rect 11564 10854 11578 10906
rect 11602 10854 11616 10906
rect 11616 10854 11628 10906
rect 11628 10854 11658 10906
rect 11682 10854 11692 10906
rect 11692 10854 11738 10906
rect 11442 10852 11498 10854
rect 11522 10852 11578 10854
rect 11602 10852 11658 10854
rect 11682 10852 11738 10854
rect 4328 10362 4384 10364
rect 4408 10362 4464 10364
rect 4488 10362 4544 10364
rect 4568 10362 4624 10364
rect 4328 10310 4374 10362
rect 4374 10310 4384 10362
rect 4408 10310 4438 10362
rect 4438 10310 4450 10362
rect 4450 10310 4464 10362
rect 4488 10310 4502 10362
rect 4502 10310 4514 10362
rect 4514 10310 4544 10362
rect 4568 10310 4578 10362
rect 4578 10310 4624 10362
rect 4328 10308 4384 10310
rect 4408 10308 4464 10310
rect 4488 10308 4544 10310
rect 4568 10308 4624 10310
rect 12102 10362 12158 10364
rect 12182 10362 12238 10364
rect 12262 10362 12318 10364
rect 12342 10362 12398 10364
rect 12102 10310 12148 10362
rect 12148 10310 12158 10362
rect 12182 10310 12212 10362
rect 12212 10310 12224 10362
rect 12224 10310 12238 10362
rect 12262 10310 12276 10362
rect 12276 10310 12288 10362
rect 12288 10310 12318 10362
rect 12342 10310 12352 10362
rect 12352 10310 12398 10362
rect 12102 10308 12158 10310
rect 12182 10308 12238 10310
rect 12262 10308 12318 10310
rect 12342 10308 12398 10310
rect 3668 9818 3724 9820
rect 3748 9818 3804 9820
rect 3828 9818 3884 9820
rect 3908 9818 3964 9820
rect 3668 9766 3714 9818
rect 3714 9766 3724 9818
rect 3748 9766 3778 9818
rect 3778 9766 3790 9818
rect 3790 9766 3804 9818
rect 3828 9766 3842 9818
rect 3842 9766 3854 9818
rect 3854 9766 3884 9818
rect 3908 9766 3918 9818
rect 3918 9766 3964 9818
rect 3668 9764 3724 9766
rect 3748 9764 3804 9766
rect 3828 9764 3884 9766
rect 3908 9764 3964 9766
rect 11442 9818 11498 9820
rect 11522 9818 11578 9820
rect 11602 9818 11658 9820
rect 11682 9818 11738 9820
rect 11442 9766 11488 9818
rect 11488 9766 11498 9818
rect 11522 9766 11552 9818
rect 11552 9766 11564 9818
rect 11564 9766 11578 9818
rect 11602 9766 11616 9818
rect 11616 9766 11628 9818
rect 11628 9766 11658 9818
rect 11682 9766 11692 9818
rect 11692 9766 11738 9818
rect 11442 9764 11498 9766
rect 11522 9764 11578 9766
rect 11602 9764 11658 9766
rect 11682 9764 11738 9766
rect 4328 9274 4384 9276
rect 4408 9274 4464 9276
rect 4488 9274 4544 9276
rect 4568 9274 4624 9276
rect 4328 9222 4374 9274
rect 4374 9222 4384 9274
rect 4408 9222 4438 9274
rect 4438 9222 4450 9274
rect 4450 9222 4464 9274
rect 4488 9222 4502 9274
rect 4502 9222 4514 9274
rect 4514 9222 4544 9274
rect 4568 9222 4578 9274
rect 4578 9222 4624 9274
rect 4328 9220 4384 9222
rect 4408 9220 4464 9222
rect 4488 9220 4544 9222
rect 4568 9220 4624 9222
rect 12102 9274 12158 9276
rect 12182 9274 12238 9276
rect 12262 9274 12318 9276
rect 12342 9274 12398 9276
rect 12102 9222 12148 9274
rect 12148 9222 12158 9274
rect 12182 9222 12212 9274
rect 12212 9222 12224 9274
rect 12224 9222 12238 9274
rect 12262 9222 12276 9274
rect 12276 9222 12288 9274
rect 12288 9222 12318 9274
rect 12342 9222 12352 9274
rect 12352 9222 12398 9274
rect 12102 9220 12158 9222
rect 12182 9220 12238 9222
rect 12262 9220 12318 9222
rect 12342 9220 12398 9222
rect 3668 8730 3724 8732
rect 3748 8730 3804 8732
rect 3828 8730 3884 8732
rect 3908 8730 3964 8732
rect 3668 8678 3714 8730
rect 3714 8678 3724 8730
rect 3748 8678 3778 8730
rect 3778 8678 3790 8730
rect 3790 8678 3804 8730
rect 3828 8678 3842 8730
rect 3842 8678 3854 8730
rect 3854 8678 3884 8730
rect 3908 8678 3918 8730
rect 3918 8678 3964 8730
rect 3668 8676 3724 8678
rect 3748 8676 3804 8678
rect 3828 8676 3884 8678
rect 3908 8676 3964 8678
rect 11442 8730 11498 8732
rect 11522 8730 11578 8732
rect 11602 8730 11658 8732
rect 11682 8730 11738 8732
rect 11442 8678 11488 8730
rect 11488 8678 11498 8730
rect 11522 8678 11552 8730
rect 11552 8678 11564 8730
rect 11564 8678 11578 8730
rect 11602 8678 11616 8730
rect 11616 8678 11628 8730
rect 11628 8678 11658 8730
rect 11682 8678 11692 8730
rect 11692 8678 11738 8730
rect 11442 8676 11498 8678
rect 11522 8676 11578 8678
rect 11602 8676 11658 8678
rect 11682 8676 11738 8678
rect 4328 8186 4384 8188
rect 4408 8186 4464 8188
rect 4488 8186 4544 8188
rect 4568 8186 4624 8188
rect 4328 8134 4374 8186
rect 4374 8134 4384 8186
rect 4408 8134 4438 8186
rect 4438 8134 4450 8186
rect 4450 8134 4464 8186
rect 4488 8134 4502 8186
rect 4502 8134 4514 8186
rect 4514 8134 4544 8186
rect 4568 8134 4578 8186
rect 4578 8134 4624 8186
rect 4328 8132 4384 8134
rect 4408 8132 4464 8134
rect 4488 8132 4544 8134
rect 4568 8132 4624 8134
rect 12102 8186 12158 8188
rect 12182 8186 12238 8188
rect 12262 8186 12318 8188
rect 12342 8186 12398 8188
rect 12102 8134 12148 8186
rect 12148 8134 12158 8186
rect 12182 8134 12212 8186
rect 12212 8134 12224 8186
rect 12224 8134 12238 8186
rect 12262 8134 12276 8186
rect 12276 8134 12288 8186
rect 12288 8134 12318 8186
rect 12342 8134 12352 8186
rect 12352 8134 12398 8186
rect 12102 8132 12158 8134
rect 12182 8132 12238 8134
rect 12262 8132 12318 8134
rect 12342 8132 12398 8134
rect 3668 7642 3724 7644
rect 3748 7642 3804 7644
rect 3828 7642 3884 7644
rect 3908 7642 3964 7644
rect 3668 7590 3714 7642
rect 3714 7590 3724 7642
rect 3748 7590 3778 7642
rect 3778 7590 3790 7642
rect 3790 7590 3804 7642
rect 3828 7590 3842 7642
rect 3842 7590 3854 7642
rect 3854 7590 3884 7642
rect 3908 7590 3918 7642
rect 3918 7590 3964 7642
rect 3668 7588 3724 7590
rect 3748 7588 3804 7590
rect 3828 7588 3884 7590
rect 3908 7588 3964 7590
rect 11442 7642 11498 7644
rect 11522 7642 11578 7644
rect 11602 7642 11658 7644
rect 11682 7642 11738 7644
rect 11442 7590 11488 7642
rect 11488 7590 11498 7642
rect 11522 7590 11552 7642
rect 11552 7590 11564 7642
rect 11564 7590 11578 7642
rect 11602 7590 11616 7642
rect 11616 7590 11628 7642
rect 11628 7590 11658 7642
rect 11682 7590 11692 7642
rect 11692 7590 11738 7642
rect 11442 7588 11498 7590
rect 11522 7588 11578 7590
rect 11602 7588 11658 7590
rect 11682 7588 11738 7590
rect 4328 7098 4384 7100
rect 4408 7098 4464 7100
rect 4488 7098 4544 7100
rect 4568 7098 4624 7100
rect 4328 7046 4374 7098
rect 4374 7046 4384 7098
rect 4408 7046 4438 7098
rect 4438 7046 4450 7098
rect 4450 7046 4464 7098
rect 4488 7046 4502 7098
rect 4502 7046 4514 7098
rect 4514 7046 4544 7098
rect 4568 7046 4578 7098
rect 4578 7046 4624 7098
rect 4328 7044 4384 7046
rect 4408 7044 4464 7046
rect 4488 7044 4544 7046
rect 4568 7044 4624 7046
rect 12102 7098 12158 7100
rect 12182 7098 12238 7100
rect 12262 7098 12318 7100
rect 12342 7098 12398 7100
rect 12102 7046 12148 7098
rect 12148 7046 12158 7098
rect 12182 7046 12212 7098
rect 12212 7046 12224 7098
rect 12224 7046 12238 7098
rect 12262 7046 12276 7098
rect 12276 7046 12288 7098
rect 12288 7046 12318 7098
rect 12342 7046 12352 7098
rect 12352 7046 12398 7098
rect 12102 7044 12158 7046
rect 12182 7044 12238 7046
rect 12262 7044 12318 7046
rect 12342 7044 12398 7046
rect 3668 6554 3724 6556
rect 3748 6554 3804 6556
rect 3828 6554 3884 6556
rect 3908 6554 3964 6556
rect 3668 6502 3714 6554
rect 3714 6502 3724 6554
rect 3748 6502 3778 6554
rect 3778 6502 3790 6554
rect 3790 6502 3804 6554
rect 3828 6502 3842 6554
rect 3842 6502 3854 6554
rect 3854 6502 3884 6554
rect 3908 6502 3918 6554
rect 3918 6502 3964 6554
rect 3668 6500 3724 6502
rect 3748 6500 3804 6502
rect 3828 6500 3884 6502
rect 3908 6500 3964 6502
rect 11442 6554 11498 6556
rect 11522 6554 11578 6556
rect 11602 6554 11658 6556
rect 11682 6554 11738 6556
rect 11442 6502 11488 6554
rect 11488 6502 11498 6554
rect 11522 6502 11552 6554
rect 11552 6502 11564 6554
rect 11564 6502 11578 6554
rect 11602 6502 11616 6554
rect 11616 6502 11628 6554
rect 11628 6502 11658 6554
rect 11682 6502 11692 6554
rect 11692 6502 11738 6554
rect 11442 6500 11498 6502
rect 11522 6500 11578 6502
rect 11602 6500 11658 6502
rect 11682 6500 11738 6502
rect 4328 6010 4384 6012
rect 4408 6010 4464 6012
rect 4488 6010 4544 6012
rect 4568 6010 4624 6012
rect 4328 5958 4374 6010
rect 4374 5958 4384 6010
rect 4408 5958 4438 6010
rect 4438 5958 4450 6010
rect 4450 5958 4464 6010
rect 4488 5958 4502 6010
rect 4502 5958 4514 6010
rect 4514 5958 4544 6010
rect 4568 5958 4578 6010
rect 4578 5958 4624 6010
rect 4328 5956 4384 5958
rect 4408 5956 4464 5958
rect 4488 5956 4544 5958
rect 4568 5956 4624 5958
rect 12102 6010 12158 6012
rect 12182 6010 12238 6012
rect 12262 6010 12318 6012
rect 12342 6010 12398 6012
rect 12102 5958 12148 6010
rect 12148 5958 12158 6010
rect 12182 5958 12212 6010
rect 12212 5958 12224 6010
rect 12224 5958 12238 6010
rect 12262 5958 12276 6010
rect 12276 5958 12288 6010
rect 12288 5958 12318 6010
rect 12342 5958 12352 6010
rect 12352 5958 12398 6010
rect 12102 5956 12158 5958
rect 12182 5956 12238 5958
rect 12262 5956 12318 5958
rect 12342 5956 12398 5958
rect 3668 5466 3724 5468
rect 3748 5466 3804 5468
rect 3828 5466 3884 5468
rect 3908 5466 3964 5468
rect 3668 5414 3714 5466
rect 3714 5414 3724 5466
rect 3748 5414 3778 5466
rect 3778 5414 3790 5466
rect 3790 5414 3804 5466
rect 3828 5414 3842 5466
rect 3842 5414 3854 5466
rect 3854 5414 3884 5466
rect 3908 5414 3918 5466
rect 3918 5414 3964 5466
rect 3668 5412 3724 5414
rect 3748 5412 3804 5414
rect 3828 5412 3884 5414
rect 3908 5412 3964 5414
rect 11442 5466 11498 5468
rect 11522 5466 11578 5468
rect 11602 5466 11658 5468
rect 11682 5466 11738 5468
rect 11442 5414 11488 5466
rect 11488 5414 11498 5466
rect 11522 5414 11552 5466
rect 11552 5414 11564 5466
rect 11564 5414 11578 5466
rect 11602 5414 11616 5466
rect 11616 5414 11628 5466
rect 11628 5414 11658 5466
rect 11682 5414 11692 5466
rect 11692 5414 11738 5466
rect 11442 5412 11498 5414
rect 11522 5412 11578 5414
rect 11602 5412 11658 5414
rect 11682 5412 11738 5414
rect 4328 4922 4384 4924
rect 4408 4922 4464 4924
rect 4488 4922 4544 4924
rect 4568 4922 4624 4924
rect 4328 4870 4374 4922
rect 4374 4870 4384 4922
rect 4408 4870 4438 4922
rect 4438 4870 4450 4922
rect 4450 4870 4464 4922
rect 4488 4870 4502 4922
rect 4502 4870 4514 4922
rect 4514 4870 4544 4922
rect 4568 4870 4578 4922
rect 4578 4870 4624 4922
rect 4328 4868 4384 4870
rect 4408 4868 4464 4870
rect 4488 4868 4544 4870
rect 4568 4868 4624 4870
rect 12102 4922 12158 4924
rect 12182 4922 12238 4924
rect 12262 4922 12318 4924
rect 12342 4922 12398 4924
rect 12102 4870 12148 4922
rect 12148 4870 12158 4922
rect 12182 4870 12212 4922
rect 12212 4870 12224 4922
rect 12224 4870 12238 4922
rect 12262 4870 12276 4922
rect 12276 4870 12288 4922
rect 12288 4870 12318 4922
rect 12342 4870 12352 4922
rect 12352 4870 12398 4922
rect 12102 4868 12158 4870
rect 12182 4868 12238 4870
rect 12262 4868 12318 4870
rect 12342 4868 12398 4870
rect 3668 4378 3724 4380
rect 3748 4378 3804 4380
rect 3828 4378 3884 4380
rect 3908 4378 3964 4380
rect 3668 4326 3714 4378
rect 3714 4326 3724 4378
rect 3748 4326 3778 4378
rect 3778 4326 3790 4378
rect 3790 4326 3804 4378
rect 3828 4326 3842 4378
rect 3842 4326 3854 4378
rect 3854 4326 3884 4378
rect 3908 4326 3918 4378
rect 3918 4326 3964 4378
rect 3668 4324 3724 4326
rect 3748 4324 3804 4326
rect 3828 4324 3884 4326
rect 3908 4324 3964 4326
rect 11442 4378 11498 4380
rect 11522 4378 11578 4380
rect 11602 4378 11658 4380
rect 11682 4378 11738 4380
rect 11442 4326 11488 4378
rect 11488 4326 11498 4378
rect 11522 4326 11552 4378
rect 11552 4326 11564 4378
rect 11564 4326 11578 4378
rect 11602 4326 11616 4378
rect 11616 4326 11628 4378
rect 11628 4326 11658 4378
rect 11682 4326 11692 4378
rect 11692 4326 11738 4378
rect 11442 4324 11498 4326
rect 11522 4324 11578 4326
rect 11602 4324 11658 4326
rect 11682 4324 11738 4326
rect 4328 3834 4384 3836
rect 4408 3834 4464 3836
rect 4488 3834 4544 3836
rect 4568 3834 4624 3836
rect 4328 3782 4374 3834
rect 4374 3782 4384 3834
rect 4408 3782 4438 3834
rect 4438 3782 4450 3834
rect 4450 3782 4464 3834
rect 4488 3782 4502 3834
rect 4502 3782 4514 3834
rect 4514 3782 4544 3834
rect 4568 3782 4578 3834
rect 4578 3782 4624 3834
rect 4328 3780 4384 3782
rect 4408 3780 4464 3782
rect 4488 3780 4544 3782
rect 4568 3780 4624 3782
rect 12102 3834 12158 3836
rect 12182 3834 12238 3836
rect 12262 3834 12318 3836
rect 12342 3834 12398 3836
rect 12102 3782 12148 3834
rect 12148 3782 12158 3834
rect 12182 3782 12212 3834
rect 12212 3782 12224 3834
rect 12224 3782 12238 3834
rect 12262 3782 12276 3834
rect 12276 3782 12288 3834
rect 12288 3782 12318 3834
rect 12342 3782 12352 3834
rect 12352 3782 12398 3834
rect 12102 3780 12158 3782
rect 12182 3780 12238 3782
rect 12262 3780 12318 3782
rect 12342 3780 12398 3782
rect 3668 3290 3724 3292
rect 3748 3290 3804 3292
rect 3828 3290 3884 3292
rect 3908 3290 3964 3292
rect 3668 3238 3714 3290
rect 3714 3238 3724 3290
rect 3748 3238 3778 3290
rect 3778 3238 3790 3290
rect 3790 3238 3804 3290
rect 3828 3238 3842 3290
rect 3842 3238 3854 3290
rect 3854 3238 3884 3290
rect 3908 3238 3918 3290
rect 3918 3238 3964 3290
rect 3668 3236 3724 3238
rect 3748 3236 3804 3238
rect 3828 3236 3884 3238
rect 3908 3236 3964 3238
rect 11442 3290 11498 3292
rect 11522 3290 11578 3292
rect 11602 3290 11658 3292
rect 11682 3290 11738 3292
rect 11442 3238 11488 3290
rect 11488 3238 11498 3290
rect 11522 3238 11552 3290
rect 11552 3238 11564 3290
rect 11564 3238 11578 3290
rect 11602 3238 11616 3290
rect 11616 3238 11628 3290
rect 11628 3238 11658 3290
rect 11682 3238 11692 3290
rect 11692 3238 11738 3290
rect 11442 3236 11498 3238
rect 11522 3236 11578 3238
rect 11602 3236 11658 3238
rect 11682 3236 11738 3238
rect 4328 2746 4384 2748
rect 4408 2746 4464 2748
rect 4488 2746 4544 2748
rect 4568 2746 4624 2748
rect 4328 2694 4374 2746
rect 4374 2694 4384 2746
rect 4408 2694 4438 2746
rect 4438 2694 4450 2746
rect 4450 2694 4464 2746
rect 4488 2694 4502 2746
rect 4502 2694 4514 2746
rect 4514 2694 4544 2746
rect 4568 2694 4578 2746
rect 4578 2694 4624 2746
rect 4328 2692 4384 2694
rect 4408 2692 4464 2694
rect 4488 2692 4544 2694
rect 4568 2692 4624 2694
rect 12102 2746 12158 2748
rect 12182 2746 12238 2748
rect 12262 2746 12318 2748
rect 12342 2746 12398 2748
rect 12102 2694 12148 2746
rect 12148 2694 12158 2746
rect 12182 2694 12212 2746
rect 12212 2694 12224 2746
rect 12224 2694 12238 2746
rect 12262 2694 12276 2746
rect 12276 2694 12288 2746
rect 12288 2694 12318 2746
rect 12342 2694 12352 2746
rect 12352 2694 12398 2746
rect 12102 2692 12158 2694
rect 12182 2692 12238 2694
rect 12262 2692 12318 2694
rect 12342 2692 12398 2694
rect 3668 2202 3724 2204
rect 3748 2202 3804 2204
rect 3828 2202 3884 2204
rect 3908 2202 3964 2204
rect 3668 2150 3714 2202
rect 3714 2150 3724 2202
rect 3748 2150 3778 2202
rect 3778 2150 3790 2202
rect 3790 2150 3804 2202
rect 3828 2150 3842 2202
rect 3842 2150 3854 2202
rect 3854 2150 3884 2202
rect 3908 2150 3918 2202
rect 3918 2150 3964 2202
rect 3668 2148 3724 2150
rect 3748 2148 3804 2150
rect 3828 2148 3884 2150
rect 3908 2148 3964 2150
rect 11442 2202 11498 2204
rect 11522 2202 11578 2204
rect 11602 2202 11658 2204
rect 11682 2202 11738 2204
rect 11442 2150 11488 2202
rect 11488 2150 11498 2202
rect 11522 2150 11552 2202
rect 11552 2150 11564 2202
rect 11564 2150 11578 2202
rect 11602 2150 11616 2202
rect 11616 2150 11628 2202
rect 11628 2150 11658 2202
rect 11682 2150 11692 2202
rect 11692 2150 11738 2202
rect 11442 2148 11498 2150
rect 11522 2148 11578 2150
rect 11602 2148 11658 2150
rect 11682 2148 11738 2150
rect 4328 1658 4384 1660
rect 4408 1658 4464 1660
rect 4488 1658 4544 1660
rect 4568 1658 4624 1660
rect 4328 1606 4374 1658
rect 4374 1606 4384 1658
rect 4408 1606 4438 1658
rect 4438 1606 4450 1658
rect 4450 1606 4464 1658
rect 4488 1606 4502 1658
rect 4502 1606 4514 1658
rect 4514 1606 4544 1658
rect 4568 1606 4578 1658
rect 4578 1606 4624 1658
rect 4328 1604 4384 1606
rect 4408 1604 4464 1606
rect 4488 1604 4544 1606
rect 4568 1604 4624 1606
rect 12102 1658 12158 1660
rect 12182 1658 12238 1660
rect 12262 1658 12318 1660
rect 12342 1658 12398 1660
rect 12102 1606 12148 1658
rect 12148 1606 12158 1658
rect 12182 1606 12212 1658
rect 12212 1606 12224 1658
rect 12224 1606 12238 1658
rect 12262 1606 12276 1658
rect 12276 1606 12288 1658
rect 12288 1606 12318 1658
rect 12342 1606 12352 1658
rect 12352 1606 12398 1658
rect 12102 1604 12158 1606
rect 12182 1604 12238 1606
rect 12262 1604 12318 1606
rect 12342 1604 12398 1606
rect 3668 1114 3724 1116
rect 3748 1114 3804 1116
rect 3828 1114 3884 1116
rect 3908 1114 3964 1116
rect 3668 1062 3714 1114
rect 3714 1062 3724 1114
rect 3748 1062 3778 1114
rect 3778 1062 3790 1114
rect 3790 1062 3804 1114
rect 3828 1062 3842 1114
rect 3842 1062 3854 1114
rect 3854 1062 3884 1114
rect 3908 1062 3918 1114
rect 3918 1062 3964 1114
rect 3668 1060 3724 1062
rect 3748 1060 3804 1062
rect 3828 1060 3884 1062
rect 3908 1060 3964 1062
rect 11442 1114 11498 1116
rect 11522 1114 11578 1116
rect 11602 1114 11658 1116
rect 11682 1114 11738 1116
rect 11442 1062 11488 1114
rect 11488 1062 11498 1114
rect 11522 1062 11552 1114
rect 11552 1062 11564 1114
rect 11564 1062 11578 1114
rect 11602 1062 11616 1114
rect 11616 1062 11628 1114
rect 11628 1062 11658 1114
rect 11682 1062 11692 1114
rect 11692 1062 11738 1114
rect 11442 1060 11498 1062
rect 11522 1060 11578 1062
rect 11602 1060 11658 1062
rect 11682 1060 11738 1062
rect 19216 17434 19272 17436
rect 19296 17434 19352 17436
rect 19376 17434 19432 17436
rect 19456 17434 19512 17436
rect 19216 17382 19262 17434
rect 19262 17382 19272 17434
rect 19296 17382 19326 17434
rect 19326 17382 19338 17434
rect 19338 17382 19352 17434
rect 19376 17382 19390 17434
rect 19390 17382 19402 17434
rect 19402 17382 19432 17434
rect 19456 17382 19466 17434
rect 19466 17382 19512 17434
rect 19216 17380 19272 17382
rect 19296 17380 19352 17382
rect 19376 17380 19432 17382
rect 19456 17380 19512 17382
rect 26990 17434 27046 17436
rect 27070 17434 27126 17436
rect 27150 17434 27206 17436
rect 27230 17434 27286 17436
rect 26990 17382 27036 17434
rect 27036 17382 27046 17434
rect 27070 17382 27100 17434
rect 27100 17382 27112 17434
rect 27112 17382 27126 17434
rect 27150 17382 27164 17434
rect 27164 17382 27176 17434
rect 27176 17382 27206 17434
rect 27230 17382 27240 17434
rect 27240 17382 27286 17434
rect 26990 17380 27046 17382
rect 27070 17380 27126 17382
rect 27150 17380 27206 17382
rect 27230 17380 27286 17382
rect 19876 16890 19932 16892
rect 19956 16890 20012 16892
rect 20036 16890 20092 16892
rect 20116 16890 20172 16892
rect 19876 16838 19922 16890
rect 19922 16838 19932 16890
rect 19956 16838 19986 16890
rect 19986 16838 19998 16890
rect 19998 16838 20012 16890
rect 20036 16838 20050 16890
rect 20050 16838 20062 16890
rect 20062 16838 20092 16890
rect 20116 16838 20126 16890
rect 20126 16838 20172 16890
rect 19876 16836 19932 16838
rect 19956 16836 20012 16838
rect 20036 16836 20092 16838
rect 20116 16836 20172 16838
rect 27650 16890 27706 16892
rect 27730 16890 27786 16892
rect 27810 16890 27866 16892
rect 27890 16890 27946 16892
rect 27650 16838 27696 16890
rect 27696 16838 27706 16890
rect 27730 16838 27760 16890
rect 27760 16838 27772 16890
rect 27772 16838 27786 16890
rect 27810 16838 27824 16890
rect 27824 16838 27836 16890
rect 27836 16838 27866 16890
rect 27890 16838 27900 16890
rect 27900 16838 27946 16890
rect 27650 16836 27706 16838
rect 27730 16836 27786 16838
rect 27810 16836 27866 16838
rect 27890 16836 27946 16838
rect 19216 16346 19272 16348
rect 19296 16346 19352 16348
rect 19376 16346 19432 16348
rect 19456 16346 19512 16348
rect 19216 16294 19262 16346
rect 19262 16294 19272 16346
rect 19296 16294 19326 16346
rect 19326 16294 19338 16346
rect 19338 16294 19352 16346
rect 19376 16294 19390 16346
rect 19390 16294 19402 16346
rect 19402 16294 19432 16346
rect 19456 16294 19466 16346
rect 19466 16294 19512 16346
rect 19216 16292 19272 16294
rect 19296 16292 19352 16294
rect 19376 16292 19432 16294
rect 19456 16292 19512 16294
rect 26990 16346 27046 16348
rect 27070 16346 27126 16348
rect 27150 16346 27206 16348
rect 27230 16346 27286 16348
rect 26990 16294 27036 16346
rect 27036 16294 27046 16346
rect 27070 16294 27100 16346
rect 27100 16294 27112 16346
rect 27112 16294 27126 16346
rect 27150 16294 27164 16346
rect 27164 16294 27176 16346
rect 27176 16294 27206 16346
rect 27230 16294 27240 16346
rect 27240 16294 27286 16346
rect 26990 16292 27046 16294
rect 27070 16292 27126 16294
rect 27150 16292 27206 16294
rect 27230 16292 27286 16294
rect 19876 15802 19932 15804
rect 19956 15802 20012 15804
rect 20036 15802 20092 15804
rect 20116 15802 20172 15804
rect 19876 15750 19922 15802
rect 19922 15750 19932 15802
rect 19956 15750 19986 15802
rect 19986 15750 19998 15802
rect 19998 15750 20012 15802
rect 20036 15750 20050 15802
rect 20050 15750 20062 15802
rect 20062 15750 20092 15802
rect 20116 15750 20126 15802
rect 20126 15750 20172 15802
rect 19876 15748 19932 15750
rect 19956 15748 20012 15750
rect 20036 15748 20092 15750
rect 20116 15748 20172 15750
rect 27650 15802 27706 15804
rect 27730 15802 27786 15804
rect 27810 15802 27866 15804
rect 27890 15802 27946 15804
rect 27650 15750 27696 15802
rect 27696 15750 27706 15802
rect 27730 15750 27760 15802
rect 27760 15750 27772 15802
rect 27772 15750 27786 15802
rect 27810 15750 27824 15802
rect 27824 15750 27836 15802
rect 27836 15750 27866 15802
rect 27890 15750 27900 15802
rect 27900 15750 27946 15802
rect 27650 15748 27706 15750
rect 27730 15748 27786 15750
rect 27810 15748 27866 15750
rect 27890 15748 27946 15750
rect 19216 15258 19272 15260
rect 19296 15258 19352 15260
rect 19376 15258 19432 15260
rect 19456 15258 19512 15260
rect 19216 15206 19262 15258
rect 19262 15206 19272 15258
rect 19296 15206 19326 15258
rect 19326 15206 19338 15258
rect 19338 15206 19352 15258
rect 19376 15206 19390 15258
rect 19390 15206 19402 15258
rect 19402 15206 19432 15258
rect 19456 15206 19466 15258
rect 19466 15206 19512 15258
rect 19216 15204 19272 15206
rect 19296 15204 19352 15206
rect 19376 15204 19432 15206
rect 19456 15204 19512 15206
rect 26990 15258 27046 15260
rect 27070 15258 27126 15260
rect 27150 15258 27206 15260
rect 27230 15258 27286 15260
rect 26990 15206 27036 15258
rect 27036 15206 27046 15258
rect 27070 15206 27100 15258
rect 27100 15206 27112 15258
rect 27112 15206 27126 15258
rect 27150 15206 27164 15258
rect 27164 15206 27176 15258
rect 27176 15206 27206 15258
rect 27230 15206 27240 15258
rect 27240 15206 27286 15258
rect 26990 15204 27046 15206
rect 27070 15204 27126 15206
rect 27150 15204 27206 15206
rect 27230 15204 27286 15206
rect 19876 14714 19932 14716
rect 19956 14714 20012 14716
rect 20036 14714 20092 14716
rect 20116 14714 20172 14716
rect 19876 14662 19922 14714
rect 19922 14662 19932 14714
rect 19956 14662 19986 14714
rect 19986 14662 19998 14714
rect 19998 14662 20012 14714
rect 20036 14662 20050 14714
rect 20050 14662 20062 14714
rect 20062 14662 20092 14714
rect 20116 14662 20126 14714
rect 20126 14662 20172 14714
rect 19876 14660 19932 14662
rect 19956 14660 20012 14662
rect 20036 14660 20092 14662
rect 20116 14660 20172 14662
rect 27650 14714 27706 14716
rect 27730 14714 27786 14716
rect 27810 14714 27866 14716
rect 27890 14714 27946 14716
rect 27650 14662 27696 14714
rect 27696 14662 27706 14714
rect 27730 14662 27760 14714
rect 27760 14662 27772 14714
rect 27772 14662 27786 14714
rect 27810 14662 27824 14714
rect 27824 14662 27836 14714
rect 27836 14662 27866 14714
rect 27890 14662 27900 14714
rect 27900 14662 27946 14714
rect 27650 14660 27706 14662
rect 27730 14660 27786 14662
rect 27810 14660 27866 14662
rect 27890 14660 27946 14662
rect 31022 14340 31078 14376
rect 31022 14320 31024 14340
rect 31024 14320 31076 14340
rect 31076 14320 31078 14340
rect 19216 14170 19272 14172
rect 19296 14170 19352 14172
rect 19376 14170 19432 14172
rect 19456 14170 19512 14172
rect 19216 14118 19262 14170
rect 19262 14118 19272 14170
rect 19296 14118 19326 14170
rect 19326 14118 19338 14170
rect 19338 14118 19352 14170
rect 19376 14118 19390 14170
rect 19390 14118 19402 14170
rect 19402 14118 19432 14170
rect 19456 14118 19466 14170
rect 19466 14118 19512 14170
rect 19216 14116 19272 14118
rect 19296 14116 19352 14118
rect 19376 14116 19432 14118
rect 19456 14116 19512 14118
rect 26990 14170 27046 14172
rect 27070 14170 27126 14172
rect 27150 14170 27206 14172
rect 27230 14170 27286 14172
rect 26990 14118 27036 14170
rect 27036 14118 27046 14170
rect 27070 14118 27100 14170
rect 27100 14118 27112 14170
rect 27112 14118 27126 14170
rect 27150 14118 27164 14170
rect 27164 14118 27176 14170
rect 27176 14118 27206 14170
rect 27230 14118 27240 14170
rect 27240 14118 27286 14170
rect 26990 14116 27046 14118
rect 27070 14116 27126 14118
rect 27150 14116 27206 14118
rect 27230 14116 27286 14118
rect 19876 13626 19932 13628
rect 19956 13626 20012 13628
rect 20036 13626 20092 13628
rect 20116 13626 20172 13628
rect 19876 13574 19922 13626
rect 19922 13574 19932 13626
rect 19956 13574 19986 13626
rect 19986 13574 19998 13626
rect 19998 13574 20012 13626
rect 20036 13574 20050 13626
rect 20050 13574 20062 13626
rect 20062 13574 20092 13626
rect 20116 13574 20126 13626
rect 20126 13574 20172 13626
rect 19876 13572 19932 13574
rect 19956 13572 20012 13574
rect 20036 13572 20092 13574
rect 20116 13572 20172 13574
rect 27650 13626 27706 13628
rect 27730 13626 27786 13628
rect 27810 13626 27866 13628
rect 27890 13626 27946 13628
rect 27650 13574 27696 13626
rect 27696 13574 27706 13626
rect 27730 13574 27760 13626
rect 27760 13574 27772 13626
rect 27772 13574 27786 13626
rect 27810 13574 27824 13626
rect 27824 13574 27836 13626
rect 27836 13574 27866 13626
rect 27890 13574 27900 13626
rect 27900 13574 27946 13626
rect 27650 13572 27706 13574
rect 27730 13572 27786 13574
rect 27810 13572 27866 13574
rect 27890 13572 27946 13574
rect 19216 13082 19272 13084
rect 19296 13082 19352 13084
rect 19376 13082 19432 13084
rect 19456 13082 19512 13084
rect 19216 13030 19262 13082
rect 19262 13030 19272 13082
rect 19296 13030 19326 13082
rect 19326 13030 19338 13082
rect 19338 13030 19352 13082
rect 19376 13030 19390 13082
rect 19390 13030 19402 13082
rect 19402 13030 19432 13082
rect 19456 13030 19466 13082
rect 19466 13030 19512 13082
rect 19216 13028 19272 13030
rect 19296 13028 19352 13030
rect 19376 13028 19432 13030
rect 19456 13028 19512 13030
rect 26990 13082 27046 13084
rect 27070 13082 27126 13084
rect 27150 13082 27206 13084
rect 27230 13082 27286 13084
rect 26990 13030 27036 13082
rect 27036 13030 27046 13082
rect 27070 13030 27100 13082
rect 27100 13030 27112 13082
rect 27112 13030 27126 13082
rect 27150 13030 27164 13082
rect 27164 13030 27176 13082
rect 27176 13030 27206 13082
rect 27230 13030 27240 13082
rect 27240 13030 27286 13082
rect 26990 13028 27046 13030
rect 27070 13028 27126 13030
rect 27150 13028 27206 13030
rect 27230 13028 27286 13030
rect 19876 12538 19932 12540
rect 19956 12538 20012 12540
rect 20036 12538 20092 12540
rect 20116 12538 20172 12540
rect 19876 12486 19922 12538
rect 19922 12486 19932 12538
rect 19956 12486 19986 12538
rect 19986 12486 19998 12538
rect 19998 12486 20012 12538
rect 20036 12486 20050 12538
rect 20050 12486 20062 12538
rect 20062 12486 20092 12538
rect 20116 12486 20126 12538
rect 20126 12486 20172 12538
rect 19876 12484 19932 12486
rect 19956 12484 20012 12486
rect 20036 12484 20092 12486
rect 20116 12484 20172 12486
rect 27650 12538 27706 12540
rect 27730 12538 27786 12540
rect 27810 12538 27866 12540
rect 27890 12538 27946 12540
rect 27650 12486 27696 12538
rect 27696 12486 27706 12538
rect 27730 12486 27760 12538
rect 27760 12486 27772 12538
rect 27772 12486 27786 12538
rect 27810 12486 27824 12538
rect 27824 12486 27836 12538
rect 27836 12486 27866 12538
rect 27890 12486 27900 12538
rect 27900 12486 27946 12538
rect 27650 12484 27706 12486
rect 27730 12484 27786 12486
rect 27810 12484 27866 12486
rect 27890 12484 27946 12486
rect 19216 11994 19272 11996
rect 19296 11994 19352 11996
rect 19376 11994 19432 11996
rect 19456 11994 19512 11996
rect 19216 11942 19262 11994
rect 19262 11942 19272 11994
rect 19296 11942 19326 11994
rect 19326 11942 19338 11994
rect 19338 11942 19352 11994
rect 19376 11942 19390 11994
rect 19390 11942 19402 11994
rect 19402 11942 19432 11994
rect 19456 11942 19466 11994
rect 19466 11942 19512 11994
rect 19216 11940 19272 11942
rect 19296 11940 19352 11942
rect 19376 11940 19432 11942
rect 19456 11940 19512 11942
rect 26990 11994 27046 11996
rect 27070 11994 27126 11996
rect 27150 11994 27206 11996
rect 27230 11994 27286 11996
rect 26990 11942 27036 11994
rect 27036 11942 27046 11994
rect 27070 11942 27100 11994
rect 27100 11942 27112 11994
rect 27112 11942 27126 11994
rect 27150 11942 27164 11994
rect 27164 11942 27176 11994
rect 27176 11942 27206 11994
rect 27230 11942 27240 11994
rect 27240 11942 27286 11994
rect 26990 11940 27046 11942
rect 27070 11940 27126 11942
rect 27150 11940 27206 11942
rect 27230 11940 27286 11942
rect 19876 11450 19932 11452
rect 19956 11450 20012 11452
rect 20036 11450 20092 11452
rect 20116 11450 20172 11452
rect 19876 11398 19922 11450
rect 19922 11398 19932 11450
rect 19956 11398 19986 11450
rect 19986 11398 19998 11450
rect 19998 11398 20012 11450
rect 20036 11398 20050 11450
rect 20050 11398 20062 11450
rect 20062 11398 20092 11450
rect 20116 11398 20126 11450
rect 20126 11398 20172 11450
rect 19876 11396 19932 11398
rect 19956 11396 20012 11398
rect 20036 11396 20092 11398
rect 20116 11396 20172 11398
rect 27650 11450 27706 11452
rect 27730 11450 27786 11452
rect 27810 11450 27866 11452
rect 27890 11450 27946 11452
rect 27650 11398 27696 11450
rect 27696 11398 27706 11450
rect 27730 11398 27760 11450
rect 27760 11398 27772 11450
rect 27772 11398 27786 11450
rect 27810 11398 27824 11450
rect 27824 11398 27836 11450
rect 27836 11398 27866 11450
rect 27890 11398 27900 11450
rect 27900 11398 27946 11450
rect 27650 11396 27706 11398
rect 27730 11396 27786 11398
rect 27810 11396 27866 11398
rect 27890 11396 27946 11398
rect 19216 10906 19272 10908
rect 19296 10906 19352 10908
rect 19376 10906 19432 10908
rect 19456 10906 19512 10908
rect 19216 10854 19262 10906
rect 19262 10854 19272 10906
rect 19296 10854 19326 10906
rect 19326 10854 19338 10906
rect 19338 10854 19352 10906
rect 19376 10854 19390 10906
rect 19390 10854 19402 10906
rect 19402 10854 19432 10906
rect 19456 10854 19466 10906
rect 19466 10854 19512 10906
rect 19216 10852 19272 10854
rect 19296 10852 19352 10854
rect 19376 10852 19432 10854
rect 19456 10852 19512 10854
rect 26990 10906 27046 10908
rect 27070 10906 27126 10908
rect 27150 10906 27206 10908
rect 27230 10906 27286 10908
rect 26990 10854 27036 10906
rect 27036 10854 27046 10906
rect 27070 10854 27100 10906
rect 27100 10854 27112 10906
rect 27112 10854 27126 10906
rect 27150 10854 27164 10906
rect 27164 10854 27176 10906
rect 27176 10854 27206 10906
rect 27230 10854 27240 10906
rect 27240 10854 27286 10906
rect 26990 10852 27046 10854
rect 27070 10852 27126 10854
rect 27150 10852 27206 10854
rect 27230 10852 27286 10854
rect 19876 10362 19932 10364
rect 19956 10362 20012 10364
rect 20036 10362 20092 10364
rect 20116 10362 20172 10364
rect 19876 10310 19922 10362
rect 19922 10310 19932 10362
rect 19956 10310 19986 10362
rect 19986 10310 19998 10362
rect 19998 10310 20012 10362
rect 20036 10310 20050 10362
rect 20050 10310 20062 10362
rect 20062 10310 20092 10362
rect 20116 10310 20126 10362
rect 20126 10310 20172 10362
rect 19876 10308 19932 10310
rect 19956 10308 20012 10310
rect 20036 10308 20092 10310
rect 20116 10308 20172 10310
rect 27650 10362 27706 10364
rect 27730 10362 27786 10364
rect 27810 10362 27866 10364
rect 27890 10362 27946 10364
rect 27650 10310 27696 10362
rect 27696 10310 27706 10362
rect 27730 10310 27760 10362
rect 27760 10310 27772 10362
rect 27772 10310 27786 10362
rect 27810 10310 27824 10362
rect 27824 10310 27836 10362
rect 27836 10310 27866 10362
rect 27890 10310 27900 10362
rect 27900 10310 27946 10362
rect 27650 10308 27706 10310
rect 27730 10308 27786 10310
rect 27810 10308 27866 10310
rect 27890 10308 27946 10310
rect 19216 9818 19272 9820
rect 19296 9818 19352 9820
rect 19376 9818 19432 9820
rect 19456 9818 19512 9820
rect 19216 9766 19262 9818
rect 19262 9766 19272 9818
rect 19296 9766 19326 9818
rect 19326 9766 19338 9818
rect 19338 9766 19352 9818
rect 19376 9766 19390 9818
rect 19390 9766 19402 9818
rect 19402 9766 19432 9818
rect 19456 9766 19466 9818
rect 19466 9766 19512 9818
rect 19216 9764 19272 9766
rect 19296 9764 19352 9766
rect 19376 9764 19432 9766
rect 19456 9764 19512 9766
rect 26990 9818 27046 9820
rect 27070 9818 27126 9820
rect 27150 9818 27206 9820
rect 27230 9818 27286 9820
rect 26990 9766 27036 9818
rect 27036 9766 27046 9818
rect 27070 9766 27100 9818
rect 27100 9766 27112 9818
rect 27112 9766 27126 9818
rect 27150 9766 27164 9818
rect 27164 9766 27176 9818
rect 27176 9766 27206 9818
rect 27230 9766 27240 9818
rect 27240 9766 27286 9818
rect 26990 9764 27046 9766
rect 27070 9764 27126 9766
rect 27150 9764 27206 9766
rect 27230 9764 27286 9766
rect 19876 9274 19932 9276
rect 19956 9274 20012 9276
rect 20036 9274 20092 9276
rect 20116 9274 20172 9276
rect 19876 9222 19922 9274
rect 19922 9222 19932 9274
rect 19956 9222 19986 9274
rect 19986 9222 19998 9274
rect 19998 9222 20012 9274
rect 20036 9222 20050 9274
rect 20050 9222 20062 9274
rect 20062 9222 20092 9274
rect 20116 9222 20126 9274
rect 20126 9222 20172 9274
rect 19876 9220 19932 9222
rect 19956 9220 20012 9222
rect 20036 9220 20092 9222
rect 20116 9220 20172 9222
rect 27650 9274 27706 9276
rect 27730 9274 27786 9276
rect 27810 9274 27866 9276
rect 27890 9274 27946 9276
rect 27650 9222 27696 9274
rect 27696 9222 27706 9274
rect 27730 9222 27760 9274
rect 27760 9222 27772 9274
rect 27772 9222 27786 9274
rect 27810 9222 27824 9274
rect 27824 9222 27836 9274
rect 27836 9222 27866 9274
rect 27890 9222 27900 9274
rect 27900 9222 27946 9274
rect 27650 9220 27706 9222
rect 27730 9220 27786 9222
rect 27810 9220 27866 9222
rect 27890 9220 27946 9222
rect 19216 8730 19272 8732
rect 19296 8730 19352 8732
rect 19376 8730 19432 8732
rect 19456 8730 19512 8732
rect 19216 8678 19262 8730
rect 19262 8678 19272 8730
rect 19296 8678 19326 8730
rect 19326 8678 19338 8730
rect 19338 8678 19352 8730
rect 19376 8678 19390 8730
rect 19390 8678 19402 8730
rect 19402 8678 19432 8730
rect 19456 8678 19466 8730
rect 19466 8678 19512 8730
rect 19216 8676 19272 8678
rect 19296 8676 19352 8678
rect 19376 8676 19432 8678
rect 19456 8676 19512 8678
rect 26990 8730 27046 8732
rect 27070 8730 27126 8732
rect 27150 8730 27206 8732
rect 27230 8730 27286 8732
rect 26990 8678 27036 8730
rect 27036 8678 27046 8730
rect 27070 8678 27100 8730
rect 27100 8678 27112 8730
rect 27112 8678 27126 8730
rect 27150 8678 27164 8730
rect 27164 8678 27176 8730
rect 27176 8678 27206 8730
rect 27230 8678 27240 8730
rect 27240 8678 27286 8730
rect 26990 8676 27046 8678
rect 27070 8676 27126 8678
rect 27150 8676 27206 8678
rect 27230 8676 27286 8678
rect 19876 8186 19932 8188
rect 19956 8186 20012 8188
rect 20036 8186 20092 8188
rect 20116 8186 20172 8188
rect 19876 8134 19922 8186
rect 19922 8134 19932 8186
rect 19956 8134 19986 8186
rect 19986 8134 19998 8186
rect 19998 8134 20012 8186
rect 20036 8134 20050 8186
rect 20050 8134 20062 8186
rect 20062 8134 20092 8186
rect 20116 8134 20126 8186
rect 20126 8134 20172 8186
rect 19876 8132 19932 8134
rect 19956 8132 20012 8134
rect 20036 8132 20092 8134
rect 20116 8132 20172 8134
rect 27650 8186 27706 8188
rect 27730 8186 27786 8188
rect 27810 8186 27866 8188
rect 27890 8186 27946 8188
rect 27650 8134 27696 8186
rect 27696 8134 27706 8186
rect 27730 8134 27760 8186
rect 27760 8134 27772 8186
rect 27772 8134 27786 8186
rect 27810 8134 27824 8186
rect 27824 8134 27836 8186
rect 27836 8134 27866 8186
rect 27890 8134 27900 8186
rect 27900 8134 27946 8186
rect 27650 8132 27706 8134
rect 27730 8132 27786 8134
rect 27810 8132 27866 8134
rect 27890 8132 27946 8134
rect 19216 7642 19272 7644
rect 19296 7642 19352 7644
rect 19376 7642 19432 7644
rect 19456 7642 19512 7644
rect 19216 7590 19262 7642
rect 19262 7590 19272 7642
rect 19296 7590 19326 7642
rect 19326 7590 19338 7642
rect 19338 7590 19352 7642
rect 19376 7590 19390 7642
rect 19390 7590 19402 7642
rect 19402 7590 19432 7642
rect 19456 7590 19466 7642
rect 19466 7590 19512 7642
rect 19216 7588 19272 7590
rect 19296 7588 19352 7590
rect 19376 7588 19432 7590
rect 19456 7588 19512 7590
rect 26990 7642 27046 7644
rect 27070 7642 27126 7644
rect 27150 7642 27206 7644
rect 27230 7642 27286 7644
rect 26990 7590 27036 7642
rect 27036 7590 27046 7642
rect 27070 7590 27100 7642
rect 27100 7590 27112 7642
rect 27112 7590 27126 7642
rect 27150 7590 27164 7642
rect 27164 7590 27176 7642
rect 27176 7590 27206 7642
rect 27230 7590 27240 7642
rect 27240 7590 27286 7642
rect 26990 7588 27046 7590
rect 27070 7588 27126 7590
rect 27150 7588 27206 7590
rect 27230 7588 27286 7590
rect 19876 7098 19932 7100
rect 19956 7098 20012 7100
rect 20036 7098 20092 7100
rect 20116 7098 20172 7100
rect 19876 7046 19922 7098
rect 19922 7046 19932 7098
rect 19956 7046 19986 7098
rect 19986 7046 19998 7098
rect 19998 7046 20012 7098
rect 20036 7046 20050 7098
rect 20050 7046 20062 7098
rect 20062 7046 20092 7098
rect 20116 7046 20126 7098
rect 20126 7046 20172 7098
rect 19876 7044 19932 7046
rect 19956 7044 20012 7046
rect 20036 7044 20092 7046
rect 20116 7044 20172 7046
rect 27650 7098 27706 7100
rect 27730 7098 27786 7100
rect 27810 7098 27866 7100
rect 27890 7098 27946 7100
rect 27650 7046 27696 7098
rect 27696 7046 27706 7098
rect 27730 7046 27760 7098
rect 27760 7046 27772 7098
rect 27772 7046 27786 7098
rect 27810 7046 27824 7098
rect 27824 7046 27836 7098
rect 27836 7046 27866 7098
rect 27890 7046 27900 7098
rect 27900 7046 27946 7098
rect 27650 7044 27706 7046
rect 27730 7044 27786 7046
rect 27810 7044 27866 7046
rect 27890 7044 27946 7046
rect 19216 6554 19272 6556
rect 19296 6554 19352 6556
rect 19376 6554 19432 6556
rect 19456 6554 19512 6556
rect 19216 6502 19262 6554
rect 19262 6502 19272 6554
rect 19296 6502 19326 6554
rect 19326 6502 19338 6554
rect 19338 6502 19352 6554
rect 19376 6502 19390 6554
rect 19390 6502 19402 6554
rect 19402 6502 19432 6554
rect 19456 6502 19466 6554
rect 19466 6502 19512 6554
rect 19216 6500 19272 6502
rect 19296 6500 19352 6502
rect 19376 6500 19432 6502
rect 19456 6500 19512 6502
rect 26990 6554 27046 6556
rect 27070 6554 27126 6556
rect 27150 6554 27206 6556
rect 27230 6554 27286 6556
rect 26990 6502 27036 6554
rect 27036 6502 27046 6554
rect 27070 6502 27100 6554
rect 27100 6502 27112 6554
rect 27112 6502 27126 6554
rect 27150 6502 27164 6554
rect 27164 6502 27176 6554
rect 27176 6502 27206 6554
rect 27230 6502 27240 6554
rect 27240 6502 27286 6554
rect 26990 6500 27046 6502
rect 27070 6500 27126 6502
rect 27150 6500 27206 6502
rect 27230 6500 27286 6502
rect 19876 6010 19932 6012
rect 19956 6010 20012 6012
rect 20036 6010 20092 6012
rect 20116 6010 20172 6012
rect 19876 5958 19922 6010
rect 19922 5958 19932 6010
rect 19956 5958 19986 6010
rect 19986 5958 19998 6010
rect 19998 5958 20012 6010
rect 20036 5958 20050 6010
rect 20050 5958 20062 6010
rect 20062 5958 20092 6010
rect 20116 5958 20126 6010
rect 20126 5958 20172 6010
rect 19876 5956 19932 5958
rect 19956 5956 20012 5958
rect 20036 5956 20092 5958
rect 20116 5956 20172 5958
rect 27650 6010 27706 6012
rect 27730 6010 27786 6012
rect 27810 6010 27866 6012
rect 27890 6010 27946 6012
rect 27650 5958 27696 6010
rect 27696 5958 27706 6010
rect 27730 5958 27760 6010
rect 27760 5958 27772 6010
rect 27772 5958 27786 6010
rect 27810 5958 27824 6010
rect 27824 5958 27836 6010
rect 27836 5958 27866 6010
rect 27890 5958 27900 6010
rect 27900 5958 27946 6010
rect 27650 5956 27706 5958
rect 27730 5956 27786 5958
rect 27810 5956 27866 5958
rect 27890 5956 27946 5958
rect 19216 5466 19272 5468
rect 19296 5466 19352 5468
rect 19376 5466 19432 5468
rect 19456 5466 19512 5468
rect 19216 5414 19262 5466
rect 19262 5414 19272 5466
rect 19296 5414 19326 5466
rect 19326 5414 19338 5466
rect 19338 5414 19352 5466
rect 19376 5414 19390 5466
rect 19390 5414 19402 5466
rect 19402 5414 19432 5466
rect 19456 5414 19466 5466
rect 19466 5414 19512 5466
rect 19216 5412 19272 5414
rect 19296 5412 19352 5414
rect 19376 5412 19432 5414
rect 19456 5412 19512 5414
rect 26990 5466 27046 5468
rect 27070 5466 27126 5468
rect 27150 5466 27206 5468
rect 27230 5466 27286 5468
rect 26990 5414 27036 5466
rect 27036 5414 27046 5466
rect 27070 5414 27100 5466
rect 27100 5414 27112 5466
rect 27112 5414 27126 5466
rect 27150 5414 27164 5466
rect 27164 5414 27176 5466
rect 27176 5414 27206 5466
rect 27230 5414 27240 5466
rect 27240 5414 27286 5466
rect 26990 5412 27046 5414
rect 27070 5412 27126 5414
rect 27150 5412 27206 5414
rect 27230 5412 27286 5414
rect 19876 4922 19932 4924
rect 19956 4922 20012 4924
rect 20036 4922 20092 4924
rect 20116 4922 20172 4924
rect 19876 4870 19922 4922
rect 19922 4870 19932 4922
rect 19956 4870 19986 4922
rect 19986 4870 19998 4922
rect 19998 4870 20012 4922
rect 20036 4870 20050 4922
rect 20050 4870 20062 4922
rect 20062 4870 20092 4922
rect 20116 4870 20126 4922
rect 20126 4870 20172 4922
rect 19876 4868 19932 4870
rect 19956 4868 20012 4870
rect 20036 4868 20092 4870
rect 20116 4868 20172 4870
rect 27650 4922 27706 4924
rect 27730 4922 27786 4924
rect 27810 4922 27866 4924
rect 27890 4922 27946 4924
rect 27650 4870 27696 4922
rect 27696 4870 27706 4922
rect 27730 4870 27760 4922
rect 27760 4870 27772 4922
rect 27772 4870 27786 4922
rect 27810 4870 27824 4922
rect 27824 4870 27836 4922
rect 27836 4870 27866 4922
rect 27890 4870 27900 4922
rect 27900 4870 27946 4922
rect 27650 4868 27706 4870
rect 27730 4868 27786 4870
rect 27810 4868 27866 4870
rect 27890 4868 27946 4870
rect 19216 4378 19272 4380
rect 19296 4378 19352 4380
rect 19376 4378 19432 4380
rect 19456 4378 19512 4380
rect 19216 4326 19262 4378
rect 19262 4326 19272 4378
rect 19296 4326 19326 4378
rect 19326 4326 19338 4378
rect 19338 4326 19352 4378
rect 19376 4326 19390 4378
rect 19390 4326 19402 4378
rect 19402 4326 19432 4378
rect 19456 4326 19466 4378
rect 19466 4326 19512 4378
rect 19216 4324 19272 4326
rect 19296 4324 19352 4326
rect 19376 4324 19432 4326
rect 19456 4324 19512 4326
rect 26990 4378 27046 4380
rect 27070 4378 27126 4380
rect 27150 4378 27206 4380
rect 27230 4378 27286 4380
rect 26990 4326 27036 4378
rect 27036 4326 27046 4378
rect 27070 4326 27100 4378
rect 27100 4326 27112 4378
rect 27112 4326 27126 4378
rect 27150 4326 27164 4378
rect 27164 4326 27176 4378
rect 27176 4326 27206 4378
rect 27230 4326 27240 4378
rect 27240 4326 27286 4378
rect 26990 4324 27046 4326
rect 27070 4324 27126 4326
rect 27150 4324 27206 4326
rect 27230 4324 27286 4326
rect 19876 3834 19932 3836
rect 19956 3834 20012 3836
rect 20036 3834 20092 3836
rect 20116 3834 20172 3836
rect 19876 3782 19922 3834
rect 19922 3782 19932 3834
rect 19956 3782 19986 3834
rect 19986 3782 19998 3834
rect 19998 3782 20012 3834
rect 20036 3782 20050 3834
rect 20050 3782 20062 3834
rect 20062 3782 20092 3834
rect 20116 3782 20126 3834
rect 20126 3782 20172 3834
rect 19876 3780 19932 3782
rect 19956 3780 20012 3782
rect 20036 3780 20092 3782
rect 20116 3780 20172 3782
rect 27650 3834 27706 3836
rect 27730 3834 27786 3836
rect 27810 3834 27866 3836
rect 27890 3834 27946 3836
rect 27650 3782 27696 3834
rect 27696 3782 27706 3834
rect 27730 3782 27760 3834
rect 27760 3782 27772 3834
rect 27772 3782 27786 3834
rect 27810 3782 27824 3834
rect 27824 3782 27836 3834
rect 27836 3782 27866 3834
rect 27890 3782 27900 3834
rect 27900 3782 27946 3834
rect 27650 3780 27706 3782
rect 27730 3780 27786 3782
rect 27810 3780 27866 3782
rect 27890 3780 27946 3782
rect 19216 3290 19272 3292
rect 19296 3290 19352 3292
rect 19376 3290 19432 3292
rect 19456 3290 19512 3292
rect 19216 3238 19262 3290
rect 19262 3238 19272 3290
rect 19296 3238 19326 3290
rect 19326 3238 19338 3290
rect 19338 3238 19352 3290
rect 19376 3238 19390 3290
rect 19390 3238 19402 3290
rect 19402 3238 19432 3290
rect 19456 3238 19466 3290
rect 19466 3238 19512 3290
rect 19216 3236 19272 3238
rect 19296 3236 19352 3238
rect 19376 3236 19432 3238
rect 19456 3236 19512 3238
rect 26990 3290 27046 3292
rect 27070 3290 27126 3292
rect 27150 3290 27206 3292
rect 27230 3290 27286 3292
rect 26990 3238 27036 3290
rect 27036 3238 27046 3290
rect 27070 3238 27100 3290
rect 27100 3238 27112 3290
rect 27112 3238 27126 3290
rect 27150 3238 27164 3290
rect 27164 3238 27176 3290
rect 27176 3238 27206 3290
rect 27230 3238 27240 3290
rect 27240 3238 27286 3290
rect 26990 3236 27046 3238
rect 27070 3236 27126 3238
rect 27150 3236 27206 3238
rect 27230 3236 27286 3238
rect 19876 2746 19932 2748
rect 19956 2746 20012 2748
rect 20036 2746 20092 2748
rect 20116 2746 20172 2748
rect 19876 2694 19922 2746
rect 19922 2694 19932 2746
rect 19956 2694 19986 2746
rect 19986 2694 19998 2746
rect 19998 2694 20012 2746
rect 20036 2694 20050 2746
rect 20050 2694 20062 2746
rect 20062 2694 20092 2746
rect 20116 2694 20126 2746
rect 20126 2694 20172 2746
rect 19876 2692 19932 2694
rect 19956 2692 20012 2694
rect 20036 2692 20092 2694
rect 20116 2692 20172 2694
rect 27650 2746 27706 2748
rect 27730 2746 27786 2748
rect 27810 2746 27866 2748
rect 27890 2746 27946 2748
rect 27650 2694 27696 2746
rect 27696 2694 27706 2746
rect 27730 2694 27760 2746
rect 27760 2694 27772 2746
rect 27772 2694 27786 2746
rect 27810 2694 27824 2746
rect 27824 2694 27836 2746
rect 27836 2694 27866 2746
rect 27890 2694 27900 2746
rect 27900 2694 27946 2746
rect 27650 2692 27706 2694
rect 27730 2692 27786 2694
rect 27810 2692 27866 2694
rect 27890 2692 27946 2694
rect 19216 2202 19272 2204
rect 19296 2202 19352 2204
rect 19376 2202 19432 2204
rect 19456 2202 19512 2204
rect 19216 2150 19262 2202
rect 19262 2150 19272 2202
rect 19296 2150 19326 2202
rect 19326 2150 19338 2202
rect 19338 2150 19352 2202
rect 19376 2150 19390 2202
rect 19390 2150 19402 2202
rect 19402 2150 19432 2202
rect 19456 2150 19466 2202
rect 19466 2150 19512 2202
rect 19216 2148 19272 2150
rect 19296 2148 19352 2150
rect 19376 2148 19432 2150
rect 19456 2148 19512 2150
rect 26990 2202 27046 2204
rect 27070 2202 27126 2204
rect 27150 2202 27206 2204
rect 27230 2202 27286 2204
rect 26990 2150 27036 2202
rect 27036 2150 27046 2202
rect 27070 2150 27100 2202
rect 27100 2150 27112 2202
rect 27112 2150 27126 2202
rect 27150 2150 27164 2202
rect 27164 2150 27176 2202
rect 27176 2150 27206 2202
rect 27230 2150 27240 2202
rect 27240 2150 27286 2202
rect 26990 2148 27046 2150
rect 27070 2148 27126 2150
rect 27150 2148 27206 2150
rect 27230 2148 27286 2150
rect 19876 1658 19932 1660
rect 19956 1658 20012 1660
rect 20036 1658 20092 1660
rect 20116 1658 20172 1660
rect 19876 1606 19922 1658
rect 19922 1606 19932 1658
rect 19956 1606 19986 1658
rect 19986 1606 19998 1658
rect 19998 1606 20012 1658
rect 20036 1606 20050 1658
rect 20050 1606 20062 1658
rect 20062 1606 20092 1658
rect 20116 1606 20126 1658
rect 20126 1606 20172 1658
rect 19876 1604 19932 1606
rect 19956 1604 20012 1606
rect 20036 1604 20092 1606
rect 20116 1604 20172 1606
rect 27650 1658 27706 1660
rect 27730 1658 27786 1660
rect 27810 1658 27866 1660
rect 27890 1658 27946 1660
rect 27650 1606 27696 1658
rect 27696 1606 27706 1658
rect 27730 1606 27760 1658
rect 27760 1606 27772 1658
rect 27772 1606 27786 1658
rect 27810 1606 27824 1658
rect 27824 1606 27836 1658
rect 27836 1606 27866 1658
rect 27890 1606 27900 1658
rect 27900 1606 27946 1658
rect 27650 1604 27706 1606
rect 27730 1604 27786 1606
rect 27810 1604 27866 1606
rect 27890 1604 27946 1606
rect 19216 1114 19272 1116
rect 19296 1114 19352 1116
rect 19376 1114 19432 1116
rect 19456 1114 19512 1116
rect 19216 1062 19262 1114
rect 19262 1062 19272 1114
rect 19296 1062 19326 1114
rect 19326 1062 19338 1114
rect 19338 1062 19352 1114
rect 19376 1062 19390 1114
rect 19390 1062 19402 1114
rect 19402 1062 19432 1114
rect 19456 1062 19466 1114
rect 19466 1062 19512 1114
rect 19216 1060 19272 1062
rect 19296 1060 19352 1062
rect 19376 1060 19432 1062
rect 19456 1060 19512 1062
rect 26990 1114 27046 1116
rect 27070 1114 27126 1116
rect 27150 1114 27206 1116
rect 27230 1114 27286 1116
rect 26990 1062 27036 1114
rect 27036 1062 27046 1114
rect 27070 1062 27100 1114
rect 27100 1062 27112 1114
rect 27112 1062 27126 1114
rect 27150 1062 27164 1114
rect 27164 1062 27176 1114
rect 27176 1062 27206 1114
rect 27230 1062 27240 1114
rect 27240 1062 27286 1114
rect 26990 1060 27046 1062
rect 27070 1060 27126 1062
rect 27150 1060 27206 1062
rect 27230 1060 27286 1062
rect 4328 570 4384 572
rect 4408 570 4464 572
rect 4488 570 4544 572
rect 4568 570 4624 572
rect 4328 518 4374 570
rect 4374 518 4384 570
rect 4408 518 4438 570
rect 4438 518 4450 570
rect 4450 518 4464 570
rect 4488 518 4502 570
rect 4502 518 4514 570
rect 4514 518 4544 570
rect 4568 518 4578 570
rect 4578 518 4624 570
rect 4328 516 4384 518
rect 4408 516 4464 518
rect 4488 516 4544 518
rect 4568 516 4624 518
rect 12102 570 12158 572
rect 12182 570 12238 572
rect 12262 570 12318 572
rect 12342 570 12398 572
rect 12102 518 12148 570
rect 12148 518 12158 570
rect 12182 518 12212 570
rect 12212 518 12224 570
rect 12224 518 12238 570
rect 12262 518 12276 570
rect 12276 518 12288 570
rect 12288 518 12318 570
rect 12342 518 12352 570
rect 12352 518 12398 570
rect 12102 516 12158 518
rect 12182 516 12238 518
rect 12262 516 12318 518
rect 12342 516 12398 518
rect 19876 570 19932 572
rect 19956 570 20012 572
rect 20036 570 20092 572
rect 20116 570 20172 572
rect 19876 518 19922 570
rect 19922 518 19932 570
rect 19956 518 19986 570
rect 19986 518 19998 570
rect 19998 518 20012 570
rect 20036 518 20050 570
rect 20050 518 20062 570
rect 20062 518 20092 570
rect 20116 518 20126 570
rect 20126 518 20172 570
rect 19876 516 19932 518
rect 19956 516 20012 518
rect 20036 516 20092 518
rect 20116 516 20172 518
rect 27650 570 27706 572
rect 27730 570 27786 572
rect 27810 570 27866 572
rect 27890 570 27946 572
rect 27650 518 27696 570
rect 27696 518 27706 570
rect 27730 518 27760 570
rect 27760 518 27772 570
rect 27772 518 27786 570
rect 27810 518 27824 570
rect 27824 518 27836 570
rect 27836 518 27866 570
rect 27890 518 27900 570
rect 27900 518 27946 570
rect 27650 516 27706 518
rect 27730 516 27786 518
rect 27810 516 27866 518
rect 27890 516 27946 518
<< metal3 >>
rect 4318 19072 4634 19073
rect 4318 19008 4324 19072
rect 4388 19008 4404 19072
rect 4468 19008 4484 19072
rect 4548 19008 4564 19072
rect 4628 19008 4634 19072
rect 4318 19007 4634 19008
rect 12092 19072 12408 19073
rect 12092 19008 12098 19072
rect 12162 19008 12178 19072
rect 12242 19008 12258 19072
rect 12322 19008 12338 19072
rect 12402 19008 12408 19072
rect 12092 19007 12408 19008
rect 19866 19072 20182 19073
rect 19866 19008 19872 19072
rect 19936 19008 19952 19072
rect 20016 19008 20032 19072
rect 20096 19008 20112 19072
rect 20176 19008 20182 19072
rect 19866 19007 20182 19008
rect 27640 19072 27956 19073
rect 27640 19008 27646 19072
rect 27710 19008 27726 19072
rect 27790 19008 27806 19072
rect 27870 19008 27886 19072
rect 27950 19008 27956 19072
rect 27640 19007 27956 19008
rect 3658 18528 3974 18529
rect 0 18458 400 18488
rect 3658 18464 3664 18528
rect 3728 18464 3744 18528
rect 3808 18464 3824 18528
rect 3888 18464 3904 18528
rect 3968 18464 3974 18528
rect 3658 18463 3974 18464
rect 11432 18528 11748 18529
rect 11432 18464 11438 18528
rect 11502 18464 11518 18528
rect 11582 18464 11598 18528
rect 11662 18464 11678 18528
rect 11742 18464 11748 18528
rect 11432 18463 11748 18464
rect 19206 18528 19522 18529
rect 19206 18464 19212 18528
rect 19276 18464 19292 18528
rect 19356 18464 19372 18528
rect 19436 18464 19452 18528
rect 19516 18464 19522 18528
rect 19206 18463 19522 18464
rect 26980 18528 27296 18529
rect 26980 18464 26986 18528
rect 27050 18464 27066 18528
rect 27130 18464 27146 18528
rect 27210 18464 27226 18528
rect 27290 18464 27296 18528
rect 26980 18463 27296 18464
rect 841 18458 907 18461
rect 0 18456 907 18458
rect 0 18400 846 18456
rect 902 18400 907 18456
rect 0 18398 907 18400
rect 0 18368 400 18398
rect 841 18395 907 18398
rect 4318 17984 4634 17985
rect 4318 17920 4324 17984
rect 4388 17920 4404 17984
rect 4468 17920 4484 17984
rect 4548 17920 4564 17984
rect 4628 17920 4634 17984
rect 4318 17919 4634 17920
rect 12092 17984 12408 17985
rect 12092 17920 12098 17984
rect 12162 17920 12178 17984
rect 12242 17920 12258 17984
rect 12322 17920 12338 17984
rect 12402 17920 12408 17984
rect 12092 17919 12408 17920
rect 19866 17984 20182 17985
rect 19866 17920 19872 17984
rect 19936 17920 19952 17984
rect 20016 17920 20032 17984
rect 20096 17920 20112 17984
rect 20176 17920 20182 17984
rect 19866 17919 20182 17920
rect 27640 17984 27956 17985
rect 27640 17920 27646 17984
rect 27710 17920 27726 17984
rect 27790 17920 27806 17984
rect 27870 17920 27886 17984
rect 27950 17920 27956 17984
rect 27640 17919 27956 17920
rect 14365 17778 14431 17781
rect 15009 17778 15075 17781
rect 14365 17776 15075 17778
rect 14365 17720 14370 17776
rect 14426 17720 15014 17776
rect 15070 17720 15075 17776
rect 14365 17718 15075 17720
rect 14365 17715 14431 17718
rect 15009 17715 15075 17718
rect 3658 17440 3974 17441
rect 3658 17376 3664 17440
rect 3728 17376 3744 17440
rect 3808 17376 3824 17440
rect 3888 17376 3904 17440
rect 3968 17376 3974 17440
rect 3658 17375 3974 17376
rect 11432 17440 11748 17441
rect 11432 17376 11438 17440
rect 11502 17376 11518 17440
rect 11582 17376 11598 17440
rect 11662 17376 11678 17440
rect 11742 17376 11748 17440
rect 11432 17375 11748 17376
rect 19206 17440 19522 17441
rect 19206 17376 19212 17440
rect 19276 17376 19292 17440
rect 19356 17376 19372 17440
rect 19436 17376 19452 17440
rect 19516 17376 19522 17440
rect 19206 17375 19522 17376
rect 26980 17440 27296 17441
rect 26980 17376 26986 17440
rect 27050 17376 27066 17440
rect 27130 17376 27146 17440
rect 27210 17376 27226 17440
rect 27290 17376 27296 17440
rect 26980 17375 27296 17376
rect 4318 16896 4634 16897
rect 4318 16832 4324 16896
rect 4388 16832 4404 16896
rect 4468 16832 4484 16896
rect 4548 16832 4564 16896
rect 4628 16832 4634 16896
rect 4318 16831 4634 16832
rect 12092 16896 12408 16897
rect 12092 16832 12098 16896
rect 12162 16832 12178 16896
rect 12242 16832 12258 16896
rect 12322 16832 12338 16896
rect 12402 16832 12408 16896
rect 12092 16831 12408 16832
rect 19866 16896 20182 16897
rect 19866 16832 19872 16896
rect 19936 16832 19952 16896
rect 20016 16832 20032 16896
rect 20096 16832 20112 16896
rect 20176 16832 20182 16896
rect 19866 16831 20182 16832
rect 27640 16896 27956 16897
rect 27640 16832 27646 16896
rect 27710 16832 27726 16896
rect 27790 16832 27806 16896
rect 27870 16832 27886 16896
rect 27950 16832 27956 16896
rect 27640 16831 27956 16832
rect 3658 16352 3974 16353
rect 3658 16288 3664 16352
rect 3728 16288 3744 16352
rect 3808 16288 3824 16352
rect 3888 16288 3904 16352
rect 3968 16288 3974 16352
rect 3658 16287 3974 16288
rect 11432 16352 11748 16353
rect 11432 16288 11438 16352
rect 11502 16288 11518 16352
rect 11582 16288 11598 16352
rect 11662 16288 11678 16352
rect 11742 16288 11748 16352
rect 11432 16287 11748 16288
rect 19206 16352 19522 16353
rect 19206 16288 19212 16352
rect 19276 16288 19292 16352
rect 19356 16288 19372 16352
rect 19436 16288 19452 16352
rect 19516 16288 19522 16352
rect 19206 16287 19522 16288
rect 26980 16352 27296 16353
rect 26980 16288 26986 16352
rect 27050 16288 27066 16352
rect 27130 16288 27146 16352
rect 27210 16288 27226 16352
rect 27290 16288 27296 16352
rect 26980 16287 27296 16288
rect 4318 15808 4634 15809
rect 4318 15744 4324 15808
rect 4388 15744 4404 15808
rect 4468 15744 4484 15808
rect 4548 15744 4564 15808
rect 4628 15744 4634 15808
rect 4318 15743 4634 15744
rect 12092 15808 12408 15809
rect 12092 15744 12098 15808
rect 12162 15744 12178 15808
rect 12242 15744 12258 15808
rect 12322 15744 12338 15808
rect 12402 15744 12408 15808
rect 12092 15743 12408 15744
rect 19866 15808 20182 15809
rect 19866 15744 19872 15808
rect 19936 15744 19952 15808
rect 20016 15744 20032 15808
rect 20096 15744 20112 15808
rect 20176 15744 20182 15808
rect 19866 15743 20182 15744
rect 27640 15808 27956 15809
rect 27640 15744 27646 15808
rect 27710 15744 27726 15808
rect 27790 15744 27806 15808
rect 27870 15744 27886 15808
rect 27950 15744 27956 15808
rect 27640 15743 27956 15744
rect 3658 15264 3974 15265
rect 3658 15200 3664 15264
rect 3728 15200 3744 15264
rect 3808 15200 3824 15264
rect 3888 15200 3904 15264
rect 3968 15200 3974 15264
rect 3658 15199 3974 15200
rect 11432 15264 11748 15265
rect 11432 15200 11438 15264
rect 11502 15200 11518 15264
rect 11582 15200 11598 15264
rect 11662 15200 11678 15264
rect 11742 15200 11748 15264
rect 11432 15199 11748 15200
rect 19206 15264 19522 15265
rect 19206 15200 19212 15264
rect 19276 15200 19292 15264
rect 19356 15200 19372 15264
rect 19436 15200 19452 15264
rect 19516 15200 19522 15264
rect 19206 15199 19522 15200
rect 26980 15264 27296 15265
rect 26980 15200 26986 15264
rect 27050 15200 27066 15264
rect 27130 15200 27146 15264
rect 27210 15200 27226 15264
rect 27290 15200 27296 15264
rect 26980 15199 27296 15200
rect 4318 14720 4634 14721
rect 4318 14656 4324 14720
rect 4388 14656 4404 14720
rect 4468 14656 4484 14720
rect 4548 14656 4564 14720
rect 4628 14656 4634 14720
rect 4318 14655 4634 14656
rect 12092 14720 12408 14721
rect 12092 14656 12098 14720
rect 12162 14656 12178 14720
rect 12242 14656 12258 14720
rect 12322 14656 12338 14720
rect 12402 14656 12408 14720
rect 12092 14655 12408 14656
rect 19866 14720 20182 14721
rect 19866 14656 19872 14720
rect 19936 14656 19952 14720
rect 20016 14656 20032 14720
rect 20096 14656 20112 14720
rect 20176 14656 20182 14720
rect 19866 14655 20182 14656
rect 27640 14720 27956 14721
rect 27640 14656 27646 14720
rect 27710 14656 27726 14720
rect 27790 14656 27806 14720
rect 27870 14656 27886 14720
rect 27950 14656 27956 14720
rect 27640 14655 27956 14656
rect 31017 14378 31083 14381
rect 31600 14378 32000 14408
rect 31017 14376 32000 14378
rect 31017 14320 31022 14376
rect 31078 14320 32000 14376
rect 31017 14318 32000 14320
rect 31017 14315 31083 14318
rect 31600 14288 32000 14318
rect 3658 14176 3974 14177
rect 3658 14112 3664 14176
rect 3728 14112 3744 14176
rect 3808 14112 3824 14176
rect 3888 14112 3904 14176
rect 3968 14112 3974 14176
rect 3658 14111 3974 14112
rect 11432 14176 11748 14177
rect 11432 14112 11438 14176
rect 11502 14112 11518 14176
rect 11582 14112 11598 14176
rect 11662 14112 11678 14176
rect 11742 14112 11748 14176
rect 11432 14111 11748 14112
rect 19206 14176 19522 14177
rect 19206 14112 19212 14176
rect 19276 14112 19292 14176
rect 19356 14112 19372 14176
rect 19436 14112 19452 14176
rect 19516 14112 19522 14176
rect 19206 14111 19522 14112
rect 26980 14176 27296 14177
rect 26980 14112 26986 14176
rect 27050 14112 27066 14176
rect 27130 14112 27146 14176
rect 27210 14112 27226 14176
rect 27290 14112 27296 14176
rect 26980 14111 27296 14112
rect 4318 13632 4634 13633
rect 4318 13568 4324 13632
rect 4388 13568 4404 13632
rect 4468 13568 4484 13632
rect 4548 13568 4564 13632
rect 4628 13568 4634 13632
rect 4318 13567 4634 13568
rect 12092 13632 12408 13633
rect 12092 13568 12098 13632
rect 12162 13568 12178 13632
rect 12242 13568 12258 13632
rect 12322 13568 12338 13632
rect 12402 13568 12408 13632
rect 12092 13567 12408 13568
rect 19866 13632 20182 13633
rect 19866 13568 19872 13632
rect 19936 13568 19952 13632
rect 20016 13568 20032 13632
rect 20096 13568 20112 13632
rect 20176 13568 20182 13632
rect 19866 13567 20182 13568
rect 27640 13632 27956 13633
rect 27640 13568 27646 13632
rect 27710 13568 27726 13632
rect 27790 13568 27806 13632
rect 27870 13568 27886 13632
rect 27950 13568 27956 13632
rect 27640 13567 27956 13568
rect 3658 13088 3974 13089
rect 3658 13024 3664 13088
rect 3728 13024 3744 13088
rect 3808 13024 3824 13088
rect 3888 13024 3904 13088
rect 3968 13024 3974 13088
rect 3658 13023 3974 13024
rect 11432 13088 11748 13089
rect 11432 13024 11438 13088
rect 11502 13024 11518 13088
rect 11582 13024 11598 13088
rect 11662 13024 11678 13088
rect 11742 13024 11748 13088
rect 11432 13023 11748 13024
rect 19206 13088 19522 13089
rect 19206 13024 19212 13088
rect 19276 13024 19292 13088
rect 19356 13024 19372 13088
rect 19436 13024 19452 13088
rect 19516 13024 19522 13088
rect 19206 13023 19522 13024
rect 26980 13088 27296 13089
rect 26980 13024 26986 13088
rect 27050 13024 27066 13088
rect 27130 13024 27146 13088
rect 27210 13024 27226 13088
rect 27290 13024 27296 13088
rect 26980 13023 27296 13024
rect 4318 12544 4634 12545
rect 4318 12480 4324 12544
rect 4388 12480 4404 12544
rect 4468 12480 4484 12544
rect 4548 12480 4564 12544
rect 4628 12480 4634 12544
rect 4318 12479 4634 12480
rect 12092 12544 12408 12545
rect 12092 12480 12098 12544
rect 12162 12480 12178 12544
rect 12242 12480 12258 12544
rect 12322 12480 12338 12544
rect 12402 12480 12408 12544
rect 12092 12479 12408 12480
rect 19866 12544 20182 12545
rect 19866 12480 19872 12544
rect 19936 12480 19952 12544
rect 20016 12480 20032 12544
rect 20096 12480 20112 12544
rect 20176 12480 20182 12544
rect 19866 12479 20182 12480
rect 27640 12544 27956 12545
rect 27640 12480 27646 12544
rect 27710 12480 27726 12544
rect 27790 12480 27806 12544
rect 27870 12480 27886 12544
rect 27950 12480 27956 12544
rect 27640 12479 27956 12480
rect 3658 12000 3974 12001
rect 3658 11936 3664 12000
rect 3728 11936 3744 12000
rect 3808 11936 3824 12000
rect 3888 11936 3904 12000
rect 3968 11936 3974 12000
rect 3658 11935 3974 11936
rect 11432 12000 11748 12001
rect 11432 11936 11438 12000
rect 11502 11936 11518 12000
rect 11582 11936 11598 12000
rect 11662 11936 11678 12000
rect 11742 11936 11748 12000
rect 11432 11935 11748 11936
rect 19206 12000 19522 12001
rect 19206 11936 19212 12000
rect 19276 11936 19292 12000
rect 19356 11936 19372 12000
rect 19436 11936 19452 12000
rect 19516 11936 19522 12000
rect 19206 11935 19522 11936
rect 26980 12000 27296 12001
rect 26980 11936 26986 12000
rect 27050 11936 27066 12000
rect 27130 11936 27146 12000
rect 27210 11936 27226 12000
rect 27290 11936 27296 12000
rect 26980 11935 27296 11936
rect 4318 11456 4634 11457
rect 4318 11392 4324 11456
rect 4388 11392 4404 11456
rect 4468 11392 4484 11456
rect 4548 11392 4564 11456
rect 4628 11392 4634 11456
rect 4318 11391 4634 11392
rect 12092 11456 12408 11457
rect 12092 11392 12098 11456
rect 12162 11392 12178 11456
rect 12242 11392 12258 11456
rect 12322 11392 12338 11456
rect 12402 11392 12408 11456
rect 12092 11391 12408 11392
rect 19866 11456 20182 11457
rect 19866 11392 19872 11456
rect 19936 11392 19952 11456
rect 20016 11392 20032 11456
rect 20096 11392 20112 11456
rect 20176 11392 20182 11456
rect 19866 11391 20182 11392
rect 27640 11456 27956 11457
rect 27640 11392 27646 11456
rect 27710 11392 27726 11456
rect 27790 11392 27806 11456
rect 27870 11392 27886 11456
rect 27950 11392 27956 11456
rect 27640 11391 27956 11392
rect 3658 10912 3974 10913
rect 3658 10848 3664 10912
rect 3728 10848 3744 10912
rect 3808 10848 3824 10912
rect 3888 10848 3904 10912
rect 3968 10848 3974 10912
rect 3658 10847 3974 10848
rect 11432 10912 11748 10913
rect 11432 10848 11438 10912
rect 11502 10848 11518 10912
rect 11582 10848 11598 10912
rect 11662 10848 11678 10912
rect 11742 10848 11748 10912
rect 11432 10847 11748 10848
rect 19206 10912 19522 10913
rect 19206 10848 19212 10912
rect 19276 10848 19292 10912
rect 19356 10848 19372 10912
rect 19436 10848 19452 10912
rect 19516 10848 19522 10912
rect 19206 10847 19522 10848
rect 26980 10912 27296 10913
rect 26980 10848 26986 10912
rect 27050 10848 27066 10912
rect 27130 10848 27146 10912
rect 27210 10848 27226 10912
rect 27290 10848 27296 10912
rect 26980 10847 27296 10848
rect 4318 10368 4634 10369
rect 4318 10304 4324 10368
rect 4388 10304 4404 10368
rect 4468 10304 4484 10368
rect 4548 10304 4564 10368
rect 4628 10304 4634 10368
rect 4318 10303 4634 10304
rect 12092 10368 12408 10369
rect 12092 10304 12098 10368
rect 12162 10304 12178 10368
rect 12242 10304 12258 10368
rect 12322 10304 12338 10368
rect 12402 10304 12408 10368
rect 12092 10303 12408 10304
rect 19866 10368 20182 10369
rect 19866 10304 19872 10368
rect 19936 10304 19952 10368
rect 20016 10304 20032 10368
rect 20096 10304 20112 10368
rect 20176 10304 20182 10368
rect 19866 10303 20182 10304
rect 27640 10368 27956 10369
rect 27640 10304 27646 10368
rect 27710 10304 27726 10368
rect 27790 10304 27806 10368
rect 27870 10304 27886 10368
rect 27950 10304 27956 10368
rect 27640 10303 27956 10304
rect 3658 9824 3974 9825
rect 3658 9760 3664 9824
rect 3728 9760 3744 9824
rect 3808 9760 3824 9824
rect 3888 9760 3904 9824
rect 3968 9760 3974 9824
rect 3658 9759 3974 9760
rect 11432 9824 11748 9825
rect 11432 9760 11438 9824
rect 11502 9760 11518 9824
rect 11582 9760 11598 9824
rect 11662 9760 11678 9824
rect 11742 9760 11748 9824
rect 11432 9759 11748 9760
rect 19206 9824 19522 9825
rect 19206 9760 19212 9824
rect 19276 9760 19292 9824
rect 19356 9760 19372 9824
rect 19436 9760 19452 9824
rect 19516 9760 19522 9824
rect 19206 9759 19522 9760
rect 26980 9824 27296 9825
rect 26980 9760 26986 9824
rect 27050 9760 27066 9824
rect 27130 9760 27146 9824
rect 27210 9760 27226 9824
rect 27290 9760 27296 9824
rect 26980 9759 27296 9760
rect 4318 9280 4634 9281
rect 4318 9216 4324 9280
rect 4388 9216 4404 9280
rect 4468 9216 4484 9280
rect 4548 9216 4564 9280
rect 4628 9216 4634 9280
rect 4318 9215 4634 9216
rect 12092 9280 12408 9281
rect 12092 9216 12098 9280
rect 12162 9216 12178 9280
rect 12242 9216 12258 9280
rect 12322 9216 12338 9280
rect 12402 9216 12408 9280
rect 12092 9215 12408 9216
rect 19866 9280 20182 9281
rect 19866 9216 19872 9280
rect 19936 9216 19952 9280
rect 20016 9216 20032 9280
rect 20096 9216 20112 9280
rect 20176 9216 20182 9280
rect 19866 9215 20182 9216
rect 27640 9280 27956 9281
rect 27640 9216 27646 9280
rect 27710 9216 27726 9280
rect 27790 9216 27806 9280
rect 27870 9216 27886 9280
rect 27950 9216 27956 9280
rect 27640 9215 27956 9216
rect 3658 8736 3974 8737
rect 3658 8672 3664 8736
rect 3728 8672 3744 8736
rect 3808 8672 3824 8736
rect 3888 8672 3904 8736
rect 3968 8672 3974 8736
rect 3658 8671 3974 8672
rect 11432 8736 11748 8737
rect 11432 8672 11438 8736
rect 11502 8672 11518 8736
rect 11582 8672 11598 8736
rect 11662 8672 11678 8736
rect 11742 8672 11748 8736
rect 11432 8671 11748 8672
rect 19206 8736 19522 8737
rect 19206 8672 19212 8736
rect 19276 8672 19292 8736
rect 19356 8672 19372 8736
rect 19436 8672 19452 8736
rect 19516 8672 19522 8736
rect 19206 8671 19522 8672
rect 26980 8736 27296 8737
rect 26980 8672 26986 8736
rect 27050 8672 27066 8736
rect 27130 8672 27146 8736
rect 27210 8672 27226 8736
rect 27290 8672 27296 8736
rect 26980 8671 27296 8672
rect 4318 8192 4634 8193
rect 4318 8128 4324 8192
rect 4388 8128 4404 8192
rect 4468 8128 4484 8192
rect 4548 8128 4564 8192
rect 4628 8128 4634 8192
rect 4318 8127 4634 8128
rect 12092 8192 12408 8193
rect 12092 8128 12098 8192
rect 12162 8128 12178 8192
rect 12242 8128 12258 8192
rect 12322 8128 12338 8192
rect 12402 8128 12408 8192
rect 12092 8127 12408 8128
rect 19866 8192 20182 8193
rect 19866 8128 19872 8192
rect 19936 8128 19952 8192
rect 20016 8128 20032 8192
rect 20096 8128 20112 8192
rect 20176 8128 20182 8192
rect 19866 8127 20182 8128
rect 27640 8192 27956 8193
rect 27640 8128 27646 8192
rect 27710 8128 27726 8192
rect 27790 8128 27806 8192
rect 27870 8128 27886 8192
rect 27950 8128 27956 8192
rect 27640 8127 27956 8128
rect 3658 7648 3974 7649
rect 3658 7584 3664 7648
rect 3728 7584 3744 7648
rect 3808 7584 3824 7648
rect 3888 7584 3904 7648
rect 3968 7584 3974 7648
rect 3658 7583 3974 7584
rect 11432 7648 11748 7649
rect 11432 7584 11438 7648
rect 11502 7584 11518 7648
rect 11582 7584 11598 7648
rect 11662 7584 11678 7648
rect 11742 7584 11748 7648
rect 11432 7583 11748 7584
rect 19206 7648 19522 7649
rect 19206 7584 19212 7648
rect 19276 7584 19292 7648
rect 19356 7584 19372 7648
rect 19436 7584 19452 7648
rect 19516 7584 19522 7648
rect 19206 7583 19522 7584
rect 26980 7648 27296 7649
rect 26980 7584 26986 7648
rect 27050 7584 27066 7648
rect 27130 7584 27146 7648
rect 27210 7584 27226 7648
rect 27290 7584 27296 7648
rect 26980 7583 27296 7584
rect 4318 7104 4634 7105
rect 4318 7040 4324 7104
rect 4388 7040 4404 7104
rect 4468 7040 4484 7104
rect 4548 7040 4564 7104
rect 4628 7040 4634 7104
rect 4318 7039 4634 7040
rect 12092 7104 12408 7105
rect 12092 7040 12098 7104
rect 12162 7040 12178 7104
rect 12242 7040 12258 7104
rect 12322 7040 12338 7104
rect 12402 7040 12408 7104
rect 12092 7039 12408 7040
rect 19866 7104 20182 7105
rect 19866 7040 19872 7104
rect 19936 7040 19952 7104
rect 20016 7040 20032 7104
rect 20096 7040 20112 7104
rect 20176 7040 20182 7104
rect 19866 7039 20182 7040
rect 27640 7104 27956 7105
rect 27640 7040 27646 7104
rect 27710 7040 27726 7104
rect 27790 7040 27806 7104
rect 27870 7040 27886 7104
rect 27950 7040 27956 7104
rect 27640 7039 27956 7040
rect 3658 6560 3974 6561
rect 3658 6496 3664 6560
rect 3728 6496 3744 6560
rect 3808 6496 3824 6560
rect 3888 6496 3904 6560
rect 3968 6496 3974 6560
rect 3658 6495 3974 6496
rect 11432 6560 11748 6561
rect 11432 6496 11438 6560
rect 11502 6496 11518 6560
rect 11582 6496 11598 6560
rect 11662 6496 11678 6560
rect 11742 6496 11748 6560
rect 11432 6495 11748 6496
rect 19206 6560 19522 6561
rect 19206 6496 19212 6560
rect 19276 6496 19292 6560
rect 19356 6496 19372 6560
rect 19436 6496 19452 6560
rect 19516 6496 19522 6560
rect 19206 6495 19522 6496
rect 26980 6560 27296 6561
rect 26980 6496 26986 6560
rect 27050 6496 27066 6560
rect 27130 6496 27146 6560
rect 27210 6496 27226 6560
rect 27290 6496 27296 6560
rect 26980 6495 27296 6496
rect 4318 6016 4634 6017
rect 4318 5952 4324 6016
rect 4388 5952 4404 6016
rect 4468 5952 4484 6016
rect 4548 5952 4564 6016
rect 4628 5952 4634 6016
rect 4318 5951 4634 5952
rect 12092 6016 12408 6017
rect 12092 5952 12098 6016
rect 12162 5952 12178 6016
rect 12242 5952 12258 6016
rect 12322 5952 12338 6016
rect 12402 5952 12408 6016
rect 12092 5951 12408 5952
rect 19866 6016 20182 6017
rect 19866 5952 19872 6016
rect 19936 5952 19952 6016
rect 20016 5952 20032 6016
rect 20096 5952 20112 6016
rect 20176 5952 20182 6016
rect 19866 5951 20182 5952
rect 27640 6016 27956 6017
rect 27640 5952 27646 6016
rect 27710 5952 27726 6016
rect 27790 5952 27806 6016
rect 27870 5952 27886 6016
rect 27950 5952 27956 6016
rect 27640 5951 27956 5952
rect 3658 5472 3974 5473
rect 3658 5408 3664 5472
rect 3728 5408 3744 5472
rect 3808 5408 3824 5472
rect 3888 5408 3904 5472
rect 3968 5408 3974 5472
rect 3658 5407 3974 5408
rect 11432 5472 11748 5473
rect 11432 5408 11438 5472
rect 11502 5408 11518 5472
rect 11582 5408 11598 5472
rect 11662 5408 11678 5472
rect 11742 5408 11748 5472
rect 11432 5407 11748 5408
rect 19206 5472 19522 5473
rect 19206 5408 19212 5472
rect 19276 5408 19292 5472
rect 19356 5408 19372 5472
rect 19436 5408 19452 5472
rect 19516 5408 19522 5472
rect 19206 5407 19522 5408
rect 26980 5472 27296 5473
rect 26980 5408 26986 5472
rect 27050 5408 27066 5472
rect 27130 5408 27146 5472
rect 27210 5408 27226 5472
rect 27290 5408 27296 5472
rect 26980 5407 27296 5408
rect 4318 4928 4634 4929
rect 4318 4864 4324 4928
rect 4388 4864 4404 4928
rect 4468 4864 4484 4928
rect 4548 4864 4564 4928
rect 4628 4864 4634 4928
rect 4318 4863 4634 4864
rect 12092 4928 12408 4929
rect 12092 4864 12098 4928
rect 12162 4864 12178 4928
rect 12242 4864 12258 4928
rect 12322 4864 12338 4928
rect 12402 4864 12408 4928
rect 12092 4863 12408 4864
rect 19866 4928 20182 4929
rect 19866 4864 19872 4928
rect 19936 4864 19952 4928
rect 20016 4864 20032 4928
rect 20096 4864 20112 4928
rect 20176 4864 20182 4928
rect 19866 4863 20182 4864
rect 27640 4928 27956 4929
rect 27640 4864 27646 4928
rect 27710 4864 27726 4928
rect 27790 4864 27806 4928
rect 27870 4864 27886 4928
rect 27950 4864 27956 4928
rect 27640 4863 27956 4864
rect 3658 4384 3974 4385
rect 3658 4320 3664 4384
rect 3728 4320 3744 4384
rect 3808 4320 3824 4384
rect 3888 4320 3904 4384
rect 3968 4320 3974 4384
rect 3658 4319 3974 4320
rect 11432 4384 11748 4385
rect 11432 4320 11438 4384
rect 11502 4320 11518 4384
rect 11582 4320 11598 4384
rect 11662 4320 11678 4384
rect 11742 4320 11748 4384
rect 11432 4319 11748 4320
rect 19206 4384 19522 4385
rect 19206 4320 19212 4384
rect 19276 4320 19292 4384
rect 19356 4320 19372 4384
rect 19436 4320 19452 4384
rect 19516 4320 19522 4384
rect 19206 4319 19522 4320
rect 26980 4384 27296 4385
rect 26980 4320 26986 4384
rect 27050 4320 27066 4384
rect 27130 4320 27146 4384
rect 27210 4320 27226 4384
rect 27290 4320 27296 4384
rect 26980 4319 27296 4320
rect 4318 3840 4634 3841
rect 4318 3776 4324 3840
rect 4388 3776 4404 3840
rect 4468 3776 4484 3840
rect 4548 3776 4564 3840
rect 4628 3776 4634 3840
rect 4318 3775 4634 3776
rect 12092 3840 12408 3841
rect 12092 3776 12098 3840
rect 12162 3776 12178 3840
rect 12242 3776 12258 3840
rect 12322 3776 12338 3840
rect 12402 3776 12408 3840
rect 12092 3775 12408 3776
rect 19866 3840 20182 3841
rect 19866 3776 19872 3840
rect 19936 3776 19952 3840
rect 20016 3776 20032 3840
rect 20096 3776 20112 3840
rect 20176 3776 20182 3840
rect 19866 3775 20182 3776
rect 27640 3840 27956 3841
rect 27640 3776 27646 3840
rect 27710 3776 27726 3840
rect 27790 3776 27806 3840
rect 27870 3776 27886 3840
rect 27950 3776 27956 3840
rect 27640 3775 27956 3776
rect 3658 3296 3974 3297
rect 3658 3232 3664 3296
rect 3728 3232 3744 3296
rect 3808 3232 3824 3296
rect 3888 3232 3904 3296
rect 3968 3232 3974 3296
rect 3658 3231 3974 3232
rect 11432 3296 11748 3297
rect 11432 3232 11438 3296
rect 11502 3232 11518 3296
rect 11582 3232 11598 3296
rect 11662 3232 11678 3296
rect 11742 3232 11748 3296
rect 11432 3231 11748 3232
rect 19206 3296 19522 3297
rect 19206 3232 19212 3296
rect 19276 3232 19292 3296
rect 19356 3232 19372 3296
rect 19436 3232 19452 3296
rect 19516 3232 19522 3296
rect 19206 3231 19522 3232
rect 26980 3296 27296 3297
rect 26980 3232 26986 3296
rect 27050 3232 27066 3296
rect 27130 3232 27146 3296
rect 27210 3232 27226 3296
rect 27290 3232 27296 3296
rect 26980 3231 27296 3232
rect 4318 2752 4634 2753
rect 4318 2688 4324 2752
rect 4388 2688 4404 2752
rect 4468 2688 4484 2752
rect 4548 2688 4564 2752
rect 4628 2688 4634 2752
rect 4318 2687 4634 2688
rect 12092 2752 12408 2753
rect 12092 2688 12098 2752
rect 12162 2688 12178 2752
rect 12242 2688 12258 2752
rect 12322 2688 12338 2752
rect 12402 2688 12408 2752
rect 12092 2687 12408 2688
rect 19866 2752 20182 2753
rect 19866 2688 19872 2752
rect 19936 2688 19952 2752
rect 20016 2688 20032 2752
rect 20096 2688 20112 2752
rect 20176 2688 20182 2752
rect 19866 2687 20182 2688
rect 27640 2752 27956 2753
rect 27640 2688 27646 2752
rect 27710 2688 27726 2752
rect 27790 2688 27806 2752
rect 27870 2688 27886 2752
rect 27950 2688 27956 2752
rect 27640 2687 27956 2688
rect 3658 2208 3974 2209
rect 3658 2144 3664 2208
rect 3728 2144 3744 2208
rect 3808 2144 3824 2208
rect 3888 2144 3904 2208
rect 3968 2144 3974 2208
rect 3658 2143 3974 2144
rect 11432 2208 11748 2209
rect 11432 2144 11438 2208
rect 11502 2144 11518 2208
rect 11582 2144 11598 2208
rect 11662 2144 11678 2208
rect 11742 2144 11748 2208
rect 11432 2143 11748 2144
rect 19206 2208 19522 2209
rect 19206 2144 19212 2208
rect 19276 2144 19292 2208
rect 19356 2144 19372 2208
rect 19436 2144 19452 2208
rect 19516 2144 19522 2208
rect 19206 2143 19522 2144
rect 26980 2208 27296 2209
rect 26980 2144 26986 2208
rect 27050 2144 27066 2208
rect 27130 2144 27146 2208
rect 27210 2144 27226 2208
rect 27290 2144 27296 2208
rect 26980 2143 27296 2144
rect 4318 1664 4634 1665
rect 4318 1600 4324 1664
rect 4388 1600 4404 1664
rect 4468 1600 4484 1664
rect 4548 1600 4564 1664
rect 4628 1600 4634 1664
rect 4318 1599 4634 1600
rect 12092 1664 12408 1665
rect 12092 1600 12098 1664
rect 12162 1600 12178 1664
rect 12242 1600 12258 1664
rect 12322 1600 12338 1664
rect 12402 1600 12408 1664
rect 12092 1599 12408 1600
rect 19866 1664 20182 1665
rect 19866 1600 19872 1664
rect 19936 1600 19952 1664
rect 20016 1600 20032 1664
rect 20096 1600 20112 1664
rect 20176 1600 20182 1664
rect 19866 1599 20182 1600
rect 27640 1664 27956 1665
rect 27640 1600 27646 1664
rect 27710 1600 27726 1664
rect 27790 1600 27806 1664
rect 27870 1600 27886 1664
rect 27950 1600 27956 1664
rect 27640 1599 27956 1600
rect 3658 1120 3974 1121
rect 3658 1056 3664 1120
rect 3728 1056 3744 1120
rect 3808 1056 3824 1120
rect 3888 1056 3904 1120
rect 3968 1056 3974 1120
rect 3658 1055 3974 1056
rect 11432 1120 11748 1121
rect 11432 1056 11438 1120
rect 11502 1056 11518 1120
rect 11582 1056 11598 1120
rect 11662 1056 11678 1120
rect 11742 1056 11748 1120
rect 11432 1055 11748 1056
rect 19206 1120 19522 1121
rect 19206 1056 19212 1120
rect 19276 1056 19292 1120
rect 19356 1056 19372 1120
rect 19436 1056 19452 1120
rect 19516 1056 19522 1120
rect 19206 1055 19522 1056
rect 26980 1120 27296 1121
rect 26980 1056 26986 1120
rect 27050 1056 27066 1120
rect 27130 1056 27146 1120
rect 27210 1056 27226 1120
rect 27290 1056 27296 1120
rect 26980 1055 27296 1056
rect 4318 576 4634 577
rect 4318 512 4324 576
rect 4388 512 4404 576
rect 4468 512 4484 576
rect 4548 512 4564 576
rect 4628 512 4634 576
rect 4318 511 4634 512
rect 12092 576 12408 577
rect 12092 512 12098 576
rect 12162 512 12178 576
rect 12242 512 12258 576
rect 12322 512 12338 576
rect 12402 512 12408 576
rect 12092 511 12408 512
rect 19866 576 20182 577
rect 19866 512 19872 576
rect 19936 512 19952 576
rect 20016 512 20032 576
rect 20096 512 20112 576
rect 20176 512 20182 576
rect 19866 511 20182 512
rect 27640 576 27956 577
rect 27640 512 27646 576
rect 27710 512 27726 576
rect 27790 512 27806 576
rect 27870 512 27886 576
rect 27950 512 27956 576
rect 27640 511 27956 512
<< via3 >>
rect 4324 19068 4388 19072
rect 4324 19012 4328 19068
rect 4328 19012 4384 19068
rect 4384 19012 4388 19068
rect 4324 19008 4388 19012
rect 4404 19068 4468 19072
rect 4404 19012 4408 19068
rect 4408 19012 4464 19068
rect 4464 19012 4468 19068
rect 4404 19008 4468 19012
rect 4484 19068 4548 19072
rect 4484 19012 4488 19068
rect 4488 19012 4544 19068
rect 4544 19012 4548 19068
rect 4484 19008 4548 19012
rect 4564 19068 4628 19072
rect 4564 19012 4568 19068
rect 4568 19012 4624 19068
rect 4624 19012 4628 19068
rect 4564 19008 4628 19012
rect 12098 19068 12162 19072
rect 12098 19012 12102 19068
rect 12102 19012 12158 19068
rect 12158 19012 12162 19068
rect 12098 19008 12162 19012
rect 12178 19068 12242 19072
rect 12178 19012 12182 19068
rect 12182 19012 12238 19068
rect 12238 19012 12242 19068
rect 12178 19008 12242 19012
rect 12258 19068 12322 19072
rect 12258 19012 12262 19068
rect 12262 19012 12318 19068
rect 12318 19012 12322 19068
rect 12258 19008 12322 19012
rect 12338 19068 12402 19072
rect 12338 19012 12342 19068
rect 12342 19012 12398 19068
rect 12398 19012 12402 19068
rect 12338 19008 12402 19012
rect 19872 19068 19936 19072
rect 19872 19012 19876 19068
rect 19876 19012 19932 19068
rect 19932 19012 19936 19068
rect 19872 19008 19936 19012
rect 19952 19068 20016 19072
rect 19952 19012 19956 19068
rect 19956 19012 20012 19068
rect 20012 19012 20016 19068
rect 19952 19008 20016 19012
rect 20032 19068 20096 19072
rect 20032 19012 20036 19068
rect 20036 19012 20092 19068
rect 20092 19012 20096 19068
rect 20032 19008 20096 19012
rect 20112 19068 20176 19072
rect 20112 19012 20116 19068
rect 20116 19012 20172 19068
rect 20172 19012 20176 19068
rect 20112 19008 20176 19012
rect 27646 19068 27710 19072
rect 27646 19012 27650 19068
rect 27650 19012 27706 19068
rect 27706 19012 27710 19068
rect 27646 19008 27710 19012
rect 27726 19068 27790 19072
rect 27726 19012 27730 19068
rect 27730 19012 27786 19068
rect 27786 19012 27790 19068
rect 27726 19008 27790 19012
rect 27806 19068 27870 19072
rect 27806 19012 27810 19068
rect 27810 19012 27866 19068
rect 27866 19012 27870 19068
rect 27806 19008 27870 19012
rect 27886 19068 27950 19072
rect 27886 19012 27890 19068
rect 27890 19012 27946 19068
rect 27946 19012 27950 19068
rect 27886 19008 27950 19012
rect 3664 18524 3728 18528
rect 3664 18468 3668 18524
rect 3668 18468 3724 18524
rect 3724 18468 3728 18524
rect 3664 18464 3728 18468
rect 3744 18524 3808 18528
rect 3744 18468 3748 18524
rect 3748 18468 3804 18524
rect 3804 18468 3808 18524
rect 3744 18464 3808 18468
rect 3824 18524 3888 18528
rect 3824 18468 3828 18524
rect 3828 18468 3884 18524
rect 3884 18468 3888 18524
rect 3824 18464 3888 18468
rect 3904 18524 3968 18528
rect 3904 18468 3908 18524
rect 3908 18468 3964 18524
rect 3964 18468 3968 18524
rect 3904 18464 3968 18468
rect 11438 18524 11502 18528
rect 11438 18468 11442 18524
rect 11442 18468 11498 18524
rect 11498 18468 11502 18524
rect 11438 18464 11502 18468
rect 11518 18524 11582 18528
rect 11518 18468 11522 18524
rect 11522 18468 11578 18524
rect 11578 18468 11582 18524
rect 11518 18464 11582 18468
rect 11598 18524 11662 18528
rect 11598 18468 11602 18524
rect 11602 18468 11658 18524
rect 11658 18468 11662 18524
rect 11598 18464 11662 18468
rect 11678 18524 11742 18528
rect 11678 18468 11682 18524
rect 11682 18468 11738 18524
rect 11738 18468 11742 18524
rect 11678 18464 11742 18468
rect 19212 18524 19276 18528
rect 19212 18468 19216 18524
rect 19216 18468 19272 18524
rect 19272 18468 19276 18524
rect 19212 18464 19276 18468
rect 19292 18524 19356 18528
rect 19292 18468 19296 18524
rect 19296 18468 19352 18524
rect 19352 18468 19356 18524
rect 19292 18464 19356 18468
rect 19372 18524 19436 18528
rect 19372 18468 19376 18524
rect 19376 18468 19432 18524
rect 19432 18468 19436 18524
rect 19372 18464 19436 18468
rect 19452 18524 19516 18528
rect 19452 18468 19456 18524
rect 19456 18468 19512 18524
rect 19512 18468 19516 18524
rect 19452 18464 19516 18468
rect 26986 18524 27050 18528
rect 26986 18468 26990 18524
rect 26990 18468 27046 18524
rect 27046 18468 27050 18524
rect 26986 18464 27050 18468
rect 27066 18524 27130 18528
rect 27066 18468 27070 18524
rect 27070 18468 27126 18524
rect 27126 18468 27130 18524
rect 27066 18464 27130 18468
rect 27146 18524 27210 18528
rect 27146 18468 27150 18524
rect 27150 18468 27206 18524
rect 27206 18468 27210 18524
rect 27146 18464 27210 18468
rect 27226 18524 27290 18528
rect 27226 18468 27230 18524
rect 27230 18468 27286 18524
rect 27286 18468 27290 18524
rect 27226 18464 27290 18468
rect 4324 17980 4388 17984
rect 4324 17924 4328 17980
rect 4328 17924 4384 17980
rect 4384 17924 4388 17980
rect 4324 17920 4388 17924
rect 4404 17980 4468 17984
rect 4404 17924 4408 17980
rect 4408 17924 4464 17980
rect 4464 17924 4468 17980
rect 4404 17920 4468 17924
rect 4484 17980 4548 17984
rect 4484 17924 4488 17980
rect 4488 17924 4544 17980
rect 4544 17924 4548 17980
rect 4484 17920 4548 17924
rect 4564 17980 4628 17984
rect 4564 17924 4568 17980
rect 4568 17924 4624 17980
rect 4624 17924 4628 17980
rect 4564 17920 4628 17924
rect 12098 17980 12162 17984
rect 12098 17924 12102 17980
rect 12102 17924 12158 17980
rect 12158 17924 12162 17980
rect 12098 17920 12162 17924
rect 12178 17980 12242 17984
rect 12178 17924 12182 17980
rect 12182 17924 12238 17980
rect 12238 17924 12242 17980
rect 12178 17920 12242 17924
rect 12258 17980 12322 17984
rect 12258 17924 12262 17980
rect 12262 17924 12318 17980
rect 12318 17924 12322 17980
rect 12258 17920 12322 17924
rect 12338 17980 12402 17984
rect 12338 17924 12342 17980
rect 12342 17924 12398 17980
rect 12398 17924 12402 17980
rect 12338 17920 12402 17924
rect 19872 17980 19936 17984
rect 19872 17924 19876 17980
rect 19876 17924 19932 17980
rect 19932 17924 19936 17980
rect 19872 17920 19936 17924
rect 19952 17980 20016 17984
rect 19952 17924 19956 17980
rect 19956 17924 20012 17980
rect 20012 17924 20016 17980
rect 19952 17920 20016 17924
rect 20032 17980 20096 17984
rect 20032 17924 20036 17980
rect 20036 17924 20092 17980
rect 20092 17924 20096 17980
rect 20032 17920 20096 17924
rect 20112 17980 20176 17984
rect 20112 17924 20116 17980
rect 20116 17924 20172 17980
rect 20172 17924 20176 17980
rect 20112 17920 20176 17924
rect 27646 17980 27710 17984
rect 27646 17924 27650 17980
rect 27650 17924 27706 17980
rect 27706 17924 27710 17980
rect 27646 17920 27710 17924
rect 27726 17980 27790 17984
rect 27726 17924 27730 17980
rect 27730 17924 27786 17980
rect 27786 17924 27790 17980
rect 27726 17920 27790 17924
rect 27806 17980 27870 17984
rect 27806 17924 27810 17980
rect 27810 17924 27866 17980
rect 27866 17924 27870 17980
rect 27806 17920 27870 17924
rect 27886 17980 27950 17984
rect 27886 17924 27890 17980
rect 27890 17924 27946 17980
rect 27946 17924 27950 17980
rect 27886 17920 27950 17924
rect 3664 17436 3728 17440
rect 3664 17380 3668 17436
rect 3668 17380 3724 17436
rect 3724 17380 3728 17436
rect 3664 17376 3728 17380
rect 3744 17436 3808 17440
rect 3744 17380 3748 17436
rect 3748 17380 3804 17436
rect 3804 17380 3808 17436
rect 3744 17376 3808 17380
rect 3824 17436 3888 17440
rect 3824 17380 3828 17436
rect 3828 17380 3884 17436
rect 3884 17380 3888 17436
rect 3824 17376 3888 17380
rect 3904 17436 3968 17440
rect 3904 17380 3908 17436
rect 3908 17380 3964 17436
rect 3964 17380 3968 17436
rect 3904 17376 3968 17380
rect 11438 17436 11502 17440
rect 11438 17380 11442 17436
rect 11442 17380 11498 17436
rect 11498 17380 11502 17436
rect 11438 17376 11502 17380
rect 11518 17436 11582 17440
rect 11518 17380 11522 17436
rect 11522 17380 11578 17436
rect 11578 17380 11582 17436
rect 11518 17376 11582 17380
rect 11598 17436 11662 17440
rect 11598 17380 11602 17436
rect 11602 17380 11658 17436
rect 11658 17380 11662 17436
rect 11598 17376 11662 17380
rect 11678 17436 11742 17440
rect 11678 17380 11682 17436
rect 11682 17380 11738 17436
rect 11738 17380 11742 17436
rect 11678 17376 11742 17380
rect 19212 17436 19276 17440
rect 19212 17380 19216 17436
rect 19216 17380 19272 17436
rect 19272 17380 19276 17436
rect 19212 17376 19276 17380
rect 19292 17436 19356 17440
rect 19292 17380 19296 17436
rect 19296 17380 19352 17436
rect 19352 17380 19356 17436
rect 19292 17376 19356 17380
rect 19372 17436 19436 17440
rect 19372 17380 19376 17436
rect 19376 17380 19432 17436
rect 19432 17380 19436 17436
rect 19372 17376 19436 17380
rect 19452 17436 19516 17440
rect 19452 17380 19456 17436
rect 19456 17380 19512 17436
rect 19512 17380 19516 17436
rect 19452 17376 19516 17380
rect 26986 17436 27050 17440
rect 26986 17380 26990 17436
rect 26990 17380 27046 17436
rect 27046 17380 27050 17436
rect 26986 17376 27050 17380
rect 27066 17436 27130 17440
rect 27066 17380 27070 17436
rect 27070 17380 27126 17436
rect 27126 17380 27130 17436
rect 27066 17376 27130 17380
rect 27146 17436 27210 17440
rect 27146 17380 27150 17436
rect 27150 17380 27206 17436
rect 27206 17380 27210 17436
rect 27146 17376 27210 17380
rect 27226 17436 27290 17440
rect 27226 17380 27230 17436
rect 27230 17380 27286 17436
rect 27286 17380 27290 17436
rect 27226 17376 27290 17380
rect 4324 16892 4388 16896
rect 4324 16836 4328 16892
rect 4328 16836 4384 16892
rect 4384 16836 4388 16892
rect 4324 16832 4388 16836
rect 4404 16892 4468 16896
rect 4404 16836 4408 16892
rect 4408 16836 4464 16892
rect 4464 16836 4468 16892
rect 4404 16832 4468 16836
rect 4484 16892 4548 16896
rect 4484 16836 4488 16892
rect 4488 16836 4544 16892
rect 4544 16836 4548 16892
rect 4484 16832 4548 16836
rect 4564 16892 4628 16896
rect 4564 16836 4568 16892
rect 4568 16836 4624 16892
rect 4624 16836 4628 16892
rect 4564 16832 4628 16836
rect 12098 16892 12162 16896
rect 12098 16836 12102 16892
rect 12102 16836 12158 16892
rect 12158 16836 12162 16892
rect 12098 16832 12162 16836
rect 12178 16892 12242 16896
rect 12178 16836 12182 16892
rect 12182 16836 12238 16892
rect 12238 16836 12242 16892
rect 12178 16832 12242 16836
rect 12258 16892 12322 16896
rect 12258 16836 12262 16892
rect 12262 16836 12318 16892
rect 12318 16836 12322 16892
rect 12258 16832 12322 16836
rect 12338 16892 12402 16896
rect 12338 16836 12342 16892
rect 12342 16836 12398 16892
rect 12398 16836 12402 16892
rect 12338 16832 12402 16836
rect 19872 16892 19936 16896
rect 19872 16836 19876 16892
rect 19876 16836 19932 16892
rect 19932 16836 19936 16892
rect 19872 16832 19936 16836
rect 19952 16892 20016 16896
rect 19952 16836 19956 16892
rect 19956 16836 20012 16892
rect 20012 16836 20016 16892
rect 19952 16832 20016 16836
rect 20032 16892 20096 16896
rect 20032 16836 20036 16892
rect 20036 16836 20092 16892
rect 20092 16836 20096 16892
rect 20032 16832 20096 16836
rect 20112 16892 20176 16896
rect 20112 16836 20116 16892
rect 20116 16836 20172 16892
rect 20172 16836 20176 16892
rect 20112 16832 20176 16836
rect 27646 16892 27710 16896
rect 27646 16836 27650 16892
rect 27650 16836 27706 16892
rect 27706 16836 27710 16892
rect 27646 16832 27710 16836
rect 27726 16892 27790 16896
rect 27726 16836 27730 16892
rect 27730 16836 27786 16892
rect 27786 16836 27790 16892
rect 27726 16832 27790 16836
rect 27806 16892 27870 16896
rect 27806 16836 27810 16892
rect 27810 16836 27866 16892
rect 27866 16836 27870 16892
rect 27806 16832 27870 16836
rect 27886 16892 27950 16896
rect 27886 16836 27890 16892
rect 27890 16836 27946 16892
rect 27946 16836 27950 16892
rect 27886 16832 27950 16836
rect 3664 16348 3728 16352
rect 3664 16292 3668 16348
rect 3668 16292 3724 16348
rect 3724 16292 3728 16348
rect 3664 16288 3728 16292
rect 3744 16348 3808 16352
rect 3744 16292 3748 16348
rect 3748 16292 3804 16348
rect 3804 16292 3808 16348
rect 3744 16288 3808 16292
rect 3824 16348 3888 16352
rect 3824 16292 3828 16348
rect 3828 16292 3884 16348
rect 3884 16292 3888 16348
rect 3824 16288 3888 16292
rect 3904 16348 3968 16352
rect 3904 16292 3908 16348
rect 3908 16292 3964 16348
rect 3964 16292 3968 16348
rect 3904 16288 3968 16292
rect 11438 16348 11502 16352
rect 11438 16292 11442 16348
rect 11442 16292 11498 16348
rect 11498 16292 11502 16348
rect 11438 16288 11502 16292
rect 11518 16348 11582 16352
rect 11518 16292 11522 16348
rect 11522 16292 11578 16348
rect 11578 16292 11582 16348
rect 11518 16288 11582 16292
rect 11598 16348 11662 16352
rect 11598 16292 11602 16348
rect 11602 16292 11658 16348
rect 11658 16292 11662 16348
rect 11598 16288 11662 16292
rect 11678 16348 11742 16352
rect 11678 16292 11682 16348
rect 11682 16292 11738 16348
rect 11738 16292 11742 16348
rect 11678 16288 11742 16292
rect 19212 16348 19276 16352
rect 19212 16292 19216 16348
rect 19216 16292 19272 16348
rect 19272 16292 19276 16348
rect 19212 16288 19276 16292
rect 19292 16348 19356 16352
rect 19292 16292 19296 16348
rect 19296 16292 19352 16348
rect 19352 16292 19356 16348
rect 19292 16288 19356 16292
rect 19372 16348 19436 16352
rect 19372 16292 19376 16348
rect 19376 16292 19432 16348
rect 19432 16292 19436 16348
rect 19372 16288 19436 16292
rect 19452 16348 19516 16352
rect 19452 16292 19456 16348
rect 19456 16292 19512 16348
rect 19512 16292 19516 16348
rect 19452 16288 19516 16292
rect 26986 16348 27050 16352
rect 26986 16292 26990 16348
rect 26990 16292 27046 16348
rect 27046 16292 27050 16348
rect 26986 16288 27050 16292
rect 27066 16348 27130 16352
rect 27066 16292 27070 16348
rect 27070 16292 27126 16348
rect 27126 16292 27130 16348
rect 27066 16288 27130 16292
rect 27146 16348 27210 16352
rect 27146 16292 27150 16348
rect 27150 16292 27206 16348
rect 27206 16292 27210 16348
rect 27146 16288 27210 16292
rect 27226 16348 27290 16352
rect 27226 16292 27230 16348
rect 27230 16292 27286 16348
rect 27286 16292 27290 16348
rect 27226 16288 27290 16292
rect 4324 15804 4388 15808
rect 4324 15748 4328 15804
rect 4328 15748 4384 15804
rect 4384 15748 4388 15804
rect 4324 15744 4388 15748
rect 4404 15804 4468 15808
rect 4404 15748 4408 15804
rect 4408 15748 4464 15804
rect 4464 15748 4468 15804
rect 4404 15744 4468 15748
rect 4484 15804 4548 15808
rect 4484 15748 4488 15804
rect 4488 15748 4544 15804
rect 4544 15748 4548 15804
rect 4484 15744 4548 15748
rect 4564 15804 4628 15808
rect 4564 15748 4568 15804
rect 4568 15748 4624 15804
rect 4624 15748 4628 15804
rect 4564 15744 4628 15748
rect 12098 15804 12162 15808
rect 12098 15748 12102 15804
rect 12102 15748 12158 15804
rect 12158 15748 12162 15804
rect 12098 15744 12162 15748
rect 12178 15804 12242 15808
rect 12178 15748 12182 15804
rect 12182 15748 12238 15804
rect 12238 15748 12242 15804
rect 12178 15744 12242 15748
rect 12258 15804 12322 15808
rect 12258 15748 12262 15804
rect 12262 15748 12318 15804
rect 12318 15748 12322 15804
rect 12258 15744 12322 15748
rect 12338 15804 12402 15808
rect 12338 15748 12342 15804
rect 12342 15748 12398 15804
rect 12398 15748 12402 15804
rect 12338 15744 12402 15748
rect 19872 15804 19936 15808
rect 19872 15748 19876 15804
rect 19876 15748 19932 15804
rect 19932 15748 19936 15804
rect 19872 15744 19936 15748
rect 19952 15804 20016 15808
rect 19952 15748 19956 15804
rect 19956 15748 20012 15804
rect 20012 15748 20016 15804
rect 19952 15744 20016 15748
rect 20032 15804 20096 15808
rect 20032 15748 20036 15804
rect 20036 15748 20092 15804
rect 20092 15748 20096 15804
rect 20032 15744 20096 15748
rect 20112 15804 20176 15808
rect 20112 15748 20116 15804
rect 20116 15748 20172 15804
rect 20172 15748 20176 15804
rect 20112 15744 20176 15748
rect 27646 15804 27710 15808
rect 27646 15748 27650 15804
rect 27650 15748 27706 15804
rect 27706 15748 27710 15804
rect 27646 15744 27710 15748
rect 27726 15804 27790 15808
rect 27726 15748 27730 15804
rect 27730 15748 27786 15804
rect 27786 15748 27790 15804
rect 27726 15744 27790 15748
rect 27806 15804 27870 15808
rect 27806 15748 27810 15804
rect 27810 15748 27866 15804
rect 27866 15748 27870 15804
rect 27806 15744 27870 15748
rect 27886 15804 27950 15808
rect 27886 15748 27890 15804
rect 27890 15748 27946 15804
rect 27946 15748 27950 15804
rect 27886 15744 27950 15748
rect 3664 15260 3728 15264
rect 3664 15204 3668 15260
rect 3668 15204 3724 15260
rect 3724 15204 3728 15260
rect 3664 15200 3728 15204
rect 3744 15260 3808 15264
rect 3744 15204 3748 15260
rect 3748 15204 3804 15260
rect 3804 15204 3808 15260
rect 3744 15200 3808 15204
rect 3824 15260 3888 15264
rect 3824 15204 3828 15260
rect 3828 15204 3884 15260
rect 3884 15204 3888 15260
rect 3824 15200 3888 15204
rect 3904 15260 3968 15264
rect 3904 15204 3908 15260
rect 3908 15204 3964 15260
rect 3964 15204 3968 15260
rect 3904 15200 3968 15204
rect 11438 15260 11502 15264
rect 11438 15204 11442 15260
rect 11442 15204 11498 15260
rect 11498 15204 11502 15260
rect 11438 15200 11502 15204
rect 11518 15260 11582 15264
rect 11518 15204 11522 15260
rect 11522 15204 11578 15260
rect 11578 15204 11582 15260
rect 11518 15200 11582 15204
rect 11598 15260 11662 15264
rect 11598 15204 11602 15260
rect 11602 15204 11658 15260
rect 11658 15204 11662 15260
rect 11598 15200 11662 15204
rect 11678 15260 11742 15264
rect 11678 15204 11682 15260
rect 11682 15204 11738 15260
rect 11738 15204 11742 15260
rect 11678 15200 11742 15204
rect 19212 15260 19276 15264
rect 19212 15204 19216 15260
rect 19216 15204 19272 15260
rect 19272 15204 19276 15260
rect 19212 15200 19276 15204
rect 19292 15260 19356 15264
rect 19292 15204 19296 15260
rect 19296 15204 19352 15260
rect 19352 15204 19356 15260
rect 19292 15200 19356 15204
rect 19372 15260 19436 15264
rect 19372 15204 19376 15260
rect 19376 15204 19432 15260
rect 19432 15204 19436 15260
rect 19372 15200 19436 15204
rect 19452 15260 19516 15264
rect 19452 15204 19456 15260
rect 19456 15204 19512 15260
rect 19512 15204 19516 15260
rect 19452 15200 19516 15204
rect 26986 15260 27050 15264
rect 26986 15204 26990 15260
rect 26990 15204 27046 15260
rect 27046 15204 27050 15260
rect 26986 15200 27050 15204
rect 27066 15260 27130 15264
rect 27066 15204 27070 15260
rect 27070 15204 27126 15260
rect 27126 15204 27130 15260
rect 27066 15200 27130 15204
rect 27146 15260 27210 15264
rect 27146 15204 27150 15260
rect 27150 15204 27206 15260
rect 27206 15204 27210 15260
rect 27146 15200 27210 15204
rect 27226 15260 27290 15264
rect 27226 15204 27230 15260
rect 27230 15204 27286 15260
rect 27286 15204 27290 15260
rect 27226 15200 27290 15204
rect 4324 14716 4388 14720
rect 4324 14660 4328 14716
rect 4328 14660 4384 14716
rect 4384 14660 4388 14716
rect 4324 14656 4388 14660
rect 4404 14716 4468 14720
rect 4404 14660 4408 14716
rect 4408 14660 4464 14716
rect 4464 14660 4468 14716
rect 4404 14656 4468 14660
rect 4484 14716 4548 14720
rect 4484 14660 4488 14716
rect 4488 14660 4544 14716
rect 4544 14660 4548 14716
rect 4484 14656 4548 14660
rect 4564 14716 4628 14720
rect 4564 14660 4568 14716
rect 4568 14660 4624 14716
rect 4624 14660 4628 14716
rect 4564 14656 4628 14660
rect 12098 14716 12162 14720
rect 12098 14660 12102 14716
rect 12102 14660 12158 14716
rect 12158 14660 12162 14716
rect 12098 14656 12162 14660
rect 12178 14716 12242 14720
rect 12178 14660 12182 14716
rect 12182 14660 12238 14716
rect 12238 14660 12242 14716
rect 12178 14656 12242 14660
rect 12258 14716 12322 14720
rect 12258 14660 12262 14716
rect 12262 14660 12318 14716
rect 12318 14660 12322 14716
rect 12258 14656 12322 14660
rect 12338 14716 12402 14720
rect 12338 14660 12342 14716
rect 12342 14660 12398 14716
rect 12398 14660 12402 14716
rect 12338 14656 12402 14660
rect 19872 14716 19936 14720
rect 19872 14660 19876 14716
rect 19876 14660 19932 14716
rect 19932 14660 19936 14716
rect 19872 14656 19936 14660
rect 19952 14716 20016 14720
rect 19952 14660 19956 14716
rect 19956 14660 20012 14716
rect 20012 14660 20016 14716
rect 19952 14656 20016 14660
rect 20032 14716 20096 14720
rect 20032 14660 20036 14716
rect 20036 14660 20092 14716
rect 20092 14660 20096 14716
rect 20032 14656 20096 14660
rect 20112 14716 20176 14720
rect 20112 14660 20116 14716
rect 20116 14660 20172 14716
rect 20172 14660 20176 14716
rect 20112 14656 20176 14660
rect 27646 14716 27710 14720
rect 27646 14660 27650 14716
rect 27650 14660 27706 14716
rect 27706 14660 27710 14716
rect 27646 14656 27710 14660
rect 27726 14716 27790 14720
rect 27726 14660 27730 14716
rect 27730 14660 27786 14716
rect 27786 14660 27790 14716
rect 27726 14656 27790 14660
rect 27806 14716 27870 14720
rect 27806 14660 27810 14716
rect 27810 14660 27866 14716
rect 27866 14660 27870 14716
rect 27806 14656 27870 14660
rect 27886 14716 27950 14720
rect 27886 14660 27890 14716
rect 27890 14660 27946 14716
rect 27946 14660 27950 14716
rect 27886 14656 27950 14660
rect 3664 14172 3728 14176
rect 3664 14116 3668 14172
rect 3668 14116 3724 14172
rect 3724 14116 3728 14172
rect 3664 14112 3728 14116
rect 3744 14172 3808 14176
rect 3744 14116 3748 14172
rect 3748 14116 3804 14172
rect 3804 14116 3808 14172
rect 3744 14112 3808 14116
rect 3824 14172 3888 14176
rect 3824 14116 3828 14172
rect 3828 14116 3884 14172
rect 3884 14116 3888 14172
rect 3824 14112 3888 14116
rect 3904 14172 3968 14176
rect 3904 14116 3908 14172
rect 3908 14116 3964 14172
rect 3964 14116 3968 14172
rect 3904 14112 3968 14116
rect 11438 14172 11502 14176
rect 11438 14116 11442 14172
rect 11442 14116 11498 14172
rect 11498 14116 11502 14172
rect 11438 14112 11502 14116
rect 11518 14172 11582 14176
rect 11518 14116 11522 14172
rect 11522 14116 11578 14172
rect 11578 14116 11582 14172
rect 11518 14112 11582 14116
rect 11598 14172 11662 14176
rect 11598 14116 11602 14172
rect 11602 14116 11658 14172
rect 11658 14116 11662 14172
rect 11598 14112 11662 14116
rect 11678 14172 11742 14176
rect 11678 14116 11682 14172
rect 11682 14116 11738 14172
rect 11738 14116 11742 14172
rect 11678 14112 11742 14116
rect 19212 14172 19276 14176
rect 19212 14116 19216 14172
rect 19216 14116 19272 14172
rect 19272 14116 19276 14172
rect 19212 14112 19276 14116
rect 19292 14172 19356 14176
rect 19292 14116 19296 14172
rect 19296 14116 19352 14172
rect 19352 14116 19356 14172
rect 19292 14112 19356 14116
rect 19372 14172 19436 14176
rect 19372 14116 19376 14172
rect 19376 14116 19432 14172
rect 19432 14116 19436 14172
rect 19372 14112 19436 14116
rect 19452 14172 19516 14176
rect 19452 14116 19456 14172
rect 19456 14116 19512 14172
rect 19512 14116 19516 14172
rect 19452 14112 19516 14116
rect 26986 14172 27050 14176
rect 26986 14116 26990 14172
rect 26990 14116 27046 14172
rect 27046 14116 27050 14172
rect 26986 14112 27050 14116
rect 27066 14172 27130 14176
rect 27066 14116 27070 14172
rect 27070 14116 27126 14172
rect 27126 14116 27130 14172
rect 27066 14112 27130 14116
rect 27146 14172 27210 14176
rect 27146 14116 27150 14172
rect 27150 14116 27206 14172
rect 27206 14116 27210 14172
rect 27146 14112 27210 14116
rect 27226 14172 27290 14176
rect 27226 14116 27230 14172
rect 27230 14116 27286 14172
rect 27286 14116 27290 14172
rect 27226 14112 27290 14116
rect 4324 13628 4388 13632
rect 4324 13572 4328 13628
rect 4328 13572 4384 13628
rect 4384 13572 4388 13628
rect 4324 13568 4388 13572
rect 4404 13628 4468 13632
rect 4404 13572 4408 13628
rect 4408 13572 4464 13628
rect 4464 13572 4468 13628
rect 4404 13568 4468 13572
rect 4484 13628 4548 13632
rect 4484 13572 4488 13628
rect 4488 13572 4544 13628
rect 4544 13572 4548 13628
rect 4484 13568 4548 13572
rect 4564 13628 4628 13632
rect 4564 13572 4568 13628
rect 4568 13572 4624 13628
rect 4624 13572 4628 13628
rect 4564 13568 4628 13572
rect 12098 13628 12162 13632
rect 12098 13572 12102 13628
rect 12102 13572 12158 13628
rect 12158 13572 12162 13628
rect 12098 13568 12162 13572
rect 12178 13628 12242 13632
rect 12178 13572 12182 13628
rect 12182 13572 12238 13628
rect 12238 13572 12242 13628
rect 12178 13568 12242 13572
rect 12258 13628 12322 13632
rect 12258 13572 12262 13628
rect 12262 13572 12318 13628
rect 12318 13572 12322 13628
rect 12258 13568 12322 13572
rect 12338 13628 12402 13632
rect 12338 13572 12342 13628
rect 12342 13572 12398 13628
rect 12398 13572 12402 13628
rect 12338 13568 12402 13572
rect 19872 13628 19936 13632
rect 19872 13572 19876 13628
rect 19876 13572 19932 13628
rect 19932 13572 19936 13628
rect 19872 13568 19936 13572
rect 19952 13628 20016 13632
rect 19952 13572 19956 13628
rect 19956 13572 20012 13628
rect 20012 13572 20016 13628
rect 19952 13568 20016 13572
rect 20032 13628 20096 13632
rect 20032 13572 20036 13628
rect 20036 13572 20092 13628
rect 20092 13572 20096 13628
rect 20032 13568 20096 13572
rect 20112 13628 20176 13632
rect 20112 13572 20116 13628
rect 20116 13572 20172 13628
rect 20172 13572 20176 13628
rect 20112 13568 20176 13572
rect 27646 13628 27710 13632
rect 27646 13572 27650 13628
rect 27650 13572 27706 13628
rect 27706 13572 27710 13628
rect 27646 13568 27710 13572
rect 27726 13628 27790 13632
rect 27726 13572 27730 13628
rect 27730 13572 27786 13628
rect 27786 13572 27790 13628
rect 27726 13568 27790 13572
rect 27806 13628 27870 13632
rect 27806 13572 27810 13628
rect 27810 13572 27866 13628
rect 27866 13572 27870 13628
rect 27806 13568 27870 13572
rect 27886 13628 27950 13632
rect 27886 13572 27890 13628
rect 27890 13572 27946 13628
rect 27946 13572 27950 13628
rect 27886 13568 27950 13572
rect 3664 13084 3728 13088
rect 3664 13028 3668 13084
rect 3668 13028 3724 13084
rect 3724 13028 3728 13084
rect 3664 13024 3728 13028
rect 3744 13084 3808 13088
rect 3744 13028 3748 13084
rect 3748 13028 3804 13084
rect 3804 13028 3808 13084
rect 3744 13024 3808 13028
rect 3824 13084 3888 13088
rect 3824 13028 3828 13084
rect 3828 13028 3884 13084
rect 3884 13028 3888 13084
rect 3824 13024 3888 13028
rect 3904 13084 3968 13088
rect 3904 13028 3908 13084
rect 3908 13028 3964 13084
rect 3964 13028 3968 13084
rect 3904 13024 3968 13028
rect 11438 13084 11502 13088
rect 11438 13028 11442 13084
rect 11442 13028 11498 13084
rect 11498 13028 11502 13084
rect 11438 13024 11502 13028
rect 11518 13084 11582 13088
rect 11518 13028 11522 13084
rect 11522 13028 11578 13084
rect 11578 13028 11582 13084
rect 11518 13024 11582 13028
rect 11598 13084 11662 13088
rect 11598 13028 11602 13084
rect 11602 13028 11658 13084
rect 11658 13028 11662 13084
rect 11598 13024 11662 13028
rect 11678 13084 11742 13088
rect 11678 13028 11682 13084
rect 11682 13028 11738 13084
rect 11738 13028 11742 13084
rect 11678 13024 11742 13028
rect 19212 13084 19276 13088
rect 19212 13028 19216 13084
rect 19216 13028 19272 13084
rect 19272 13028 19276 13084
rect 19212 13024 19276 13028
rect 19292 13084 19356 13088
rect 19292 13028 19296 13084
rect 19296 13028 19352 13084
rect 19352 13028 19356 13084
rect 19292 13024 19356 13028
rect 19372 13084 19436 13088
rect 19372 13028 19376 13084
rect 19376 13028 19432 13084
rect 19432 13028 19436 13084
rect 19372 13024 19436 13028
rect 19452 13084 19516 13088
rect 19452 13028 19456 13084
rect 19456 13028 19512 13084
rect 19512 13028 19516 13084
rect 19452 13024 19516 13028
rect 26986 13084 27050 13088
rect 26986 13028 26990 13084
rect 26990 13028 27046 13084
rect 27046 13028 27050 13084
rect 26986 13024 27050 13028
rect 27066 13084 27130 13088
rect 27066 13028 27070 13084
rect 27070 13028 27126 13084
rect 27126 13028 27130 13084
rect 27066 13024 27130 13028
rect 27146 13084 27210 13088
rect 27146 13028 27150 13084
rect 27150 13028 27206 13084
rect 27206 13028 27210 13084
rect 27146 13024 27210 13028
rect 27226 13084 27290 13088
rect 27226 13028 27230 13084
rect 27230 13028 27286 13084
rect 27286 13028 27290 13084
rect 27226 13024 27290 13028
rect 4324 12540 4388 12544
rect 4324 12484 4328 12540
rect 4328 12484 4384 12540
rect 4384 12484 4388 12540
rect 4324 12480 4388 12484
rect 4404 12540 4468 12544
rect 4404 12484 4408 12540
rect 4408 12484 4464 12540
rect 4464 12484 4468 12540
rect 4404 12480 4468 12484
rect 4484 12540 4548 12544
rect 4484 12484 4488 12540
rect 4488 12484 4544 12540
rect 4544 12484 4548 12540
rect 4484 12480 4548 12484
rect 4564 12540 4628 12544
rect 4564 12484 4568 12540
rect 4568 12484 4624 12540
rect 4624 12484 4628 12540
rect 4564 12480 4628 12484
rect 12098 12540 12162 12544
rect 12098 12484 12102 12540
rect 12102 12484 12158 12540
rect 12158 12484 12162 12540
rect 12098 12480 12162 12484
rect 12178 12540 12242 12544
rect 12178 12484 12182 12540
rect 12182 12484 12238 12540
rect 12238 12484 12242 12540
rect 12178 12480 12242 12484
rect 12258 12540 12322 12544
rect 12258 12484 12262 12540
rect 12262 12484 12318 12540
rect 12318 12484 12322 12540
rect 12258 12480 12322 12484
rect 12338 12540 12402 12544
rect 12338 12484 12342 12540
rect 12342 12484 12398 12540
rect 12398 12484 12402 12540
rect 12338 12480 12402 12484
rect 19872 12540 19936 12544
rect 19872 12484 19876 12540
rect 19876 12484 19932 12540
rect 19932 12484 19936 12540
rect 19872 12480 19936 12484
rect 19952 12540 20016 12544
rect 19952 12484 19956 12540
rect 19956 12484 20012 12540
rect 20012 12484 20016 12540
rect 19952 12480 20016 12484
rect 20032 12540 20096 12544
rect 20032 12484 20036 12540
rect 20036 12484 20092 12540
rect 20092 12484 20096 12540
rect 20032 12480 20096 12484
rect 20112 12540 20176 12544
rect 20112 12484 20116 12540
rect 20116 12484 20172 12540
rect 20172 12484 20176 12540
rect 20112 12480 20176 12484
rect 27646 12540 27710 12544
rect 27646 12484 27650 12540
rect 27650 12484 27706 12540
rect 27706 12484 27710 12540
rect 27646 12480 27710 12484
rect 27726 12540 27790 12544
rect 27726 12484 27730 12540
rect 27730 12484 27786 12540
rect 27786 12484 27790 12540
rect 27726 12480 27790 12484
rect 27806 12540 27870 12544
rect 27806 12484 27810 12540
rect 27810 12484 27866 12540
rect 27866 12484 27870 12540
rect 27806 12480 27870 12484
rect 27886 12540 27950 12544
rect 27886 12484 27890 12540
rect 27890 12484 27946 12540
rect 27946 12484 27950 12540
rect 27886 12480 27950 12484
rect 3664 11996 3728 12000
rect 3664 11940 3668 11996
rect 3668 11940 3724 11996
rect 3724 11940 3728 11996
rect 3664 11936 3728 11940
rect 3744 11996 3808 12000
rect 3744 11940 3748 11996
rect 3748 11940 3804 11996
rect 3804 11940 3808 11996
rect 3744 11936 3808 11940
rect 3824 11996 3888 12000
rect 3824 11940 3828 11996
rect 3828 11940 3884 11996
rect 3884 11940 3888 11996
rect 3824 11936 3888 11940
rect 3904 11996 3968 12000
rect 3904 11940 3908 11996
rect 3908 11940 3964 11996
rect 3964 11940 3968 11996
rect 3904 11936 3968 11940
rect 11438 11996 11502 12000
rect 11438 11940 11442 11996
rect 11442 11940 11498 11996
rect 11498 11940 11502 11996
rect 11438 11936 11502 11940
rect 11518 11996 11582 12000
rect 11518 11940 11522 11996
rect 11522 11940 11578 11996
rect 11578 11940 11582 11996
rect 11518 11936 11582 11940
rect 11598 11996 11662 12000
rect 11598 11940 11602 11996
rect 11602 11940 11658 11996
rect 11658 11940 11662 11996
rect 11598 11936 11662 11940
rect 11678 11996 11742 12000
rect 11678 11940 11682 11996
rect 11682 11940 11738 11996
rect 11738 11940 11742 11996
rect 11678 11936 11742 11940
rect 19212 11996 19276 12000
rect 19212 11940 19216 11996
rect 19216 11940 19272 11996
rect 19272 11940 19276 11996
rect 19212 11936 19276 11940
rect 19292 11996 19356 12000
rect 19292 11940 19296 11996
rect 19296 11940 19352 11996
rect 19352 11940 19356 11996
rect 19292 11936 19356 11940
rect 19372 11996 19436 12000
rect 19372 11940 19376 11996
rect 19376 11940 19432 11996
rect 19432 11940 19436 11996
rect 19372 11936 19436 11940
rect 19452 11996 19516 12000
rect 19452 11940 19456 11996
rect 19456 11940 19512 11996
rect 19512 11940 19516 11996
rect 19452 11936 19516 11940
rect 26986 11996 27050 12000
rect 26986 11940 26990 11996
rect 26990 11940 27046 11996
rect 27046 11940 27050 11996
rect 26986 11936 27050 11940
rect 27066 11996 27130 12000
rect 27066 11940 27070 11996
rect 27070 11940 27126 11996
rect 27126 11940 27130 11996
rect 27066 11936 27130 11940
rect 27146 11996 27210 12000
rect 27146 11940 27150 11996
rect 27150 11940 27206 11996
rect 27206 11940 27210 11996
rect 27146 11936 27210 11940
rect 27226 11996 27290 12000
rect 27226 11940 27230 11996
rect 27230 11940 27286 11996
rect 27286 11940 27290 11996
rect 27226 11936 27290 11940
rect 4324 11452 4388 11456
rect 4324 11396 4328 11452
rect 4328 11396 4384 11452
rect 4384 11396 4388 11452
rect 4324 11392 4388 11396
rect 4404 11452 4468 11456
rect 4404 11396 4408 11452
rect 4408 11396 4464 11452
rect 4464 11396 4468 11452
rect 4404 11392 4468 11396
rect 4484 11452 4548 11456
rect 4484 11396 4488 11452
rect 4488 11396 4544 11452
rect 4544 11396 4548 11452
rect 4484 11392 4548 11396
rect 4564 11452 4628 11456
rect 4564 11396 4568 11452
rect 4568 11396 4624 11452
rect 4624 11396 4628 11452
rect 4564 11392 4628 11396
rect 12098 11452 12162 11456
rect 12098 11396 12102 11452
rect 12102 11396 12158 11452
rect 12158 11396 12162 11452
rect 12098 11392 12162 11396
rect 12178 11452 12242 11456
rect 12178 11396 12182 11452
rect 12182 11396 12238 11452
rect 12238 11396 12242 11452
rect 12178 11392 12242 11396
rect 12258 11452 12322 11456
rect 12258 11396 12262 11452
rect 12262 11396 12318 11452
rect 12318 11396 12322 11452
rect 12258 11392 12322 11396
rect 12338 11452 12402 11456
rect 12338 11396 12342 11452
rect 12342 11396 12398 11452
rect 12398 11396 12402 11452
rect 12338 11392 12402 11396
rect 19872 11452 19936 11456
rect 19872 11396 19876 11452
rect 19876 11396 19932 11452
rect 19932 11396 19936 11452
rect 19872 11392 19936 11396
rect 19952 11452 20016 11456
rect 19952 11396 19956 11452
rect 19956 11396 20012 11452
rect 20012 11396 20016 11452
rect 19952 11392 20016 11396
rect 20032 11452 20096 11456
rect 20032 11396 20036 11452
rect 20036 11396 20092 11452
rect 20092 11396 20096 11452
rect 20032 11392 20096 11396
rect 20112 11452 20176 11456
rect 20112 11396 20116 11452
rect 20116 11396 20172 11452
rect 20172 11396 20176 11452
rect 20112 11392 20176 11396
rect 27646 11452 27710 11456
rect 27646 11396 27650 11452
rect 27650 11396 27706 11452
rect 27706 11396 27710 11452
rect 27646 11392 27710 11396
rect 27726 11452 27790 11456
rect 27726 11396 27730 11452
rect 27730 11396 27786 11452
rect 27786 11396 27790 11452
rect 27726 11392 27790 11396
rect 27806 11452 27870 11456
rect 27806 11396 27810 11452
rect 27810 11396 27866 11452
rect 27866 11396 27870 11452
rect 27806 11392 27870 11396
rect 27886 11452 27950 11456
rect 27886 11396 27890 11452
rect 27890 11396 27946 11452
rect 27946 11396 27950 11452
rect 27886 11392 27950 11396
rect 3664 10908 3728 10912
rect 3664 10852 3668 10908
rect 3668 10852 3724 10908
rect 3724 10852 3728 10908
rect 3664 10848 3728 10852
rect 3744 10908 3808 10912
rect 3744 10852 3748 10908
rect 3748 10852 3804 10908
rect 3804 10852 3808 10908
rect 3744 10848 3808 10852
rect 3824 10908 3888 10912
rect 3824 10852 3828 10908
rect 3828 10852 3884 10908
rect 3884 10852 3888 10908
rect 3824 10848 3888 10852
rect 3904 10908 3968 10912
rect 3904 10852 3908 10908
rect 3908 10852 3964 10908
rect 3964 10852 3968 10908
rect 3904 10848 3968 10852
rect 11438 10908 11502 10912
rect 11438 10852 11442 10908
rect 11442 10852 11498 10908
rect 11498 10852 11502 10908
rect 11438 10848 11502 10852
rect 11518 10908 11582 10912
rect 11518 10852 11522 10908
rect 11522 10852 11578 10908
rect 11578 10852 11582 10908
rect 11518 10848 11582 10852
rect 11598 10908 11662 10912
rect 11598 10852 11602 10908
rect 11602 10852 11658 10908
rect 11658 10852 11662 10908
rect 11598 10848 11662 10852
rect 11678 10908 11742 10912
rect 11678 10852 11682 10908
rect 11682 10852 11738 10908
rect 11738 10852 11742 10908
rect 11678 10848 11742 10852
rect 19212 10908 19276 10912
rect 19212 10852 19216 10908
rect 19216 10852 19272 10908
rect 19272 10852 19276 10908
rect 19212 10848 19276 10852
rect 19292 10908 19356 10912
rect 19292 10852 19296 10908
rect 19296 10852 19352 10908
rect 19352 10852 19356 10908
rect 19292 10848 19356 10852
rect 19372 10908 19436 10912
rect 19372 10852 19376 10908
rect 19376 10852 19432 10908
rect 19432 10852 19436 10908
rect 19372 10848 19436 10852
rect 19452 10908 19516 10912
rect 19452 10852 19456 10908
rect 19456 10852 19512 10908
rect 19512 10852 19516 10908
rect 19452 10848 19516 10852
rect 26986 10908 27050 10912
rect 26986 10852 26990 10908
rect 26990 10852 27046 10908
rect 27046 10852 27050 10908
rect 26986 10848 27050 10852
rect 27066 10908 27130 10912
rect 27066 10852 27070 10908
rect 27070 10852 27126 10908
rect 27126 10852 27130 10908
rect 27066 10848 27130 10852
rect 27146 10908 27210 10912
rect 27146 10852 27150 10908
rect 27150 10852 27206 10908
rect 27206 10852 27210 10908
rect 27146 10848 27210 10852
rect 27226 10908 27290 10912
rect 27226 10852 27230 10908
rect 27230 10852 27286 10908
rect 27286 10852 27290 10908
rect 27226 10848 27290 10852
rect 4324 10364 4388 10368
rect 4324 10308 4328 10364
rect 4328 10308 4384 10364
rect 4384 10308 4388 10364
rect 4324 10304 4388 10308
rect 4404 10364 4468 10368
rect 4404 10308 4408 10364
rect 4408 10308 4464 10364
rect 4464 10308 4468 10364
rect 4404 10304 4468 10308
rect 4484 10364 4548 10368
rect 4484 10308 4488 10364
rect 4488 10308 4544 10364
rect 4544 10308 4548 10364
rect 4484 10304 4548 10308
rect 4564 10364 4628 10368
rect 4564 10308 4568 10364
rect 4568 10308 4624 10364
rect 4624 10308 4628 10364
rect 4564 10304 4628 10308
rect 12098 10364 12162 10368
rect 12098 10308 12102 10364
rect 12102 10308 12158 10364
rect 12158 10308 12162 10364
rect 12098 10304 12162 10308
rect 12178 10364 12242 10368
rect 12178 10308 12182 10364
rect 12182 10308 12238 10364
rect 12238 10308 12242 10364
rect 12178 10304 12242 10308
rect 12258 10364 12322 10368
rect 12258 10308 12262 10364
rect 12262 10308 12318 10364
rect 12318 10308 12322 10364
rect 12258 10304 12322 10308
rect 12338 10364 12402 10368
rect 12338 10308 12342 10364
rect 12342 10308 12398 10364
rect 12398 10308 12402 10364
rect 12338 10304 12402 10308
rect 19872 10364 19936 10368
rect 19872 10308 19876 10364
rect 19876 10308 19932 10364
rect 19932 10308 19936 10364
rect 19872 10304 19936 10308
rect 19952 10364 20016 10368
rect 19952 10308 19956 10364
rect 19956 10308 20012 10364
rect 20012 10308 20016 10364
rect 19952 10304 20016 10308
rect 20032 10364 20096 10368
rect 20032 10308 20036 10364
rect 20036 10308 20092 10364
rect 20092 10308 20096 10364
rect 20032 10304 20096 10308
rect 20112 10364 20176 10368
rect 20112 10308 20116 10364
rect 20116 10308 20172 10364
rect 20172 10308 20176 10364
rect 20112 10304 20176 10308
rect 27646 10364 27710 10368
rect 27646 10308 27650 10364
rect 27650 10308 27706 10364
rect 27706 10308 27710 10364
rect 27646 10304 27710 10308
rect 27726 10364 27790 10368
rect 27726 10308 27730 10364
rect 27730 10308 27786 10364
rect 27786 10308 27790 10364
rect 27726 10304 27790 10308
rect 27806 10364 27870 10368
rect 27806 10308 27810 10364
rect 27810 10308 27866 10364
rect 27866 10308 27870 10364
rect 27806 10304 27870 10308
rect 27886 10364 27950 10368
rect 27886 10308 27890 10364
rect 27890 10308 27946 10364
rect 27946 10308 27950 10364
rect 27886 10304 27950 10308
rect 3664 9820 3728 9824
rect 3664 9764 3668 9820
rect 3668 9764 3724 9820
rect 3724 9764 3728 9820
rect 3664 9760 3728 9764
rect 3744 9820 3808 9824
rect 3744 9764 3748 9820
rect 3748 9764 3804 9820
rect 3804 9764 3808 9820
rect 3744 9760 3808 9764
rect 3824 9820 3888 9824
rect 3824 9764 3828 9820
rect 3828 9764 3884 9820
rect 3884 9764 3888 9820
rect 3824 9760 3888 9764
rect 3904 9820 3968 9824
rect 3904 9764 3908 9820
rect 3908 9764 3964 9820
rect 3964 9764 3968 9820
rect 3904 9760 3968 9764
rect 11438 9820 11502 9824
rect 11438 9764 11442 9820
rect 11442 9764 11498 9820
rect 11498 9764 11502 9820
rect 11438 9760 11502 9764
rect 11518 9820 11582 9824
rect 11518 9764 11522 9820
rect 11522 9764 11578 9820
rect 11578 9764 11582 9820
rect 11518 9760 11582 9764
rect 11598 9820 11662 9824
rect 11598 9764 11602 9820
rect 11602 9764 11658 9820
rect 11658 9764 11662 9820
rect 11598 9760 11662 9764
rect 11678 9820 11742 9824
rect 11678 9764 11682 9820
rect 11682 9764 11738 9820
rect 11738 9764 11742 9820
rect 11678 9760 11742 9764
rect 19212 9820 19276 9824
rect 19212 9764 19216 9820
rect 19216 9764 19272 9820
rect 19272 9764 19276 9820
rect 19212 9760 19276 9764
rect 19292 9820 19356 9824
rect 19292 9764 19296 9820
rect 19296 9764 19352 9820
rect 19352 9764 19356 9820
rect 19292 9760 19356 9764
rect 19372 9820 19436 9824
rect 19372 9764 19376 9820
rect 19376 9764 19432 9820
rect 19432 9764 19436 9820
rect 19372 9760 19436 9764
rect 19452 9820 19516 9824
rect 19452 9764 19456 9820
rect 19456 9764 19512 9820
rect 19512 9764 19516 9820
rect 19452 9760 19516 9764
rect 26986 9820 27050 9824
rect 26986 9764 26990 9820
rect 26990 9764 27046 9820
rect 27046 9764 27050 9820
rect 26986 9760 27050 9764
rect 27066 9820 27130 9824
rect 27066 9764 27070 9820
rect 27070 9764 27126 9820
rect 27126 9764 27130 9820
rect 27066 9760 27130 9764
rect 27146 9820 27210 9824
rect 27146 9764 27150 9820
rect 27150 9764 27206 9820
rect 27206 9764 27210 9820
rect 27146 9760 27210 9764
rect 27226 9820 27290 9824
rect 27226 9764 27230 9820
rect 27230 9764 27286 9820
rect 27286 9764 27290 9820
rect 27226 9760 27290 9764
rect 4324 9276 4388 9280
rect 4324 9220 4328 9276
rect 4328 9220 4384 9276
rect 4384 9220 4388 9276
rect 4324 9216 4388 9220
rect 4404 9276 4468 9280
rect 4404 9220 4408 9276
rect 4408 9220 4464 9276
rect 4464 9220 4468 9276
rect 4404 9216 4468 9220
rect 4484 9276 4548 9280
rect 4484 9220 4488 9276
rect 4488 9220 4544 9276
rect 4544 9220 4548 9276
rect 4484 9216 4548 9220
rect 4564 9276 4628 9280
rect 4564 9220 4568 9276
rect 4568 9220 4624 9276
rect 4624 9220 4628 9276
rect 4564 9216 4628 9220
rect 12098 9276 12162 9280
rect 12098 9220 12102 9276
rect 12102 9220 12158 9276
rect 12158 9220 12162 9276
rect 12098 9216 12162 9220
rect 12178 9276 12242 9280
rect 12178 9220 12182 9276
rect 12182 9220 12238 9276
rect 12238 9220 12242 9276
rect 12178 9216 12242 9220
rect 12258 9276 12322 9280
rect 12258 9220 12262 9276
rect 12262 9220 12318 9276
rect 12318 9220 12322 9276
rect 12258 9216 12322 9220
rect 12338 9276 12402 9280
rect 12338 9220 12342 9276
rect 12342 9220 12398 9276
rect 12398 9220 12402 9276
rect 12338 9216 12402 9220
rect 19872 9276 19936 9280
rect 19872 9220 19876 9276
rect 19876 9220 19932 9276
rect 19932 9220 19936 9276
rect 19872 9216 19936 9220
rect 19952 9276 20016 9280
rect 19952 9220 19956 9276
rect 19956 9220 20012 9276
rect 20012 9220 20016 9276
rect 19952 9216 20016 9220
rect 20032 9276 20096 9280
rect 20032 9220 20036 9276
rect 20036 9220 20092 9276
rect 20092 9220 20096 9276
rect 20032 9216 20096 9220
rect 20112 9276 20176 9280
rect 20112 9220 20116 9276
rect 20116 9220 20172 9276
rect 20172 9220 20176 9276
rect 20112 9216 20176 9220
rect 27646 9276 27710 9280
rect 27646 9220 27650 9276
rect 27650 9220 27706 9276
rect 27706 9220 27710 9276
rect 27646 9216 27710 9220
rect 27726 9276 27790 9280
rect 27726 9220 27730 9276
rect 27730 9220 27786 9276
rect 27786 9220 27790 9276
rect 27726 9216 27790 9220
rect 27806 9276 27870 9280
rect 27806 9220 27810 9276
rect 27810 9220 27866 9276
rect 27866 9220 27870 9276
rect 27806 9216 27870 9220
rect 27886 9276 27950 9280
rect 27886 9220 27890 9276
rect 27890 9220 27946 9276
rect 27946 9220 27950 9276
rect 27886 9216 27950 9220
rect 3664 8732 3728 8736
rect 3664 8676 3668 8732
rect 3668 8676 3724 8732
rect 3724 8676 3728 8732
rect 3664 8672 3728 8676
rect 3744 8732 3808 8736
rect 3744 8676 3748 8732
rect 3748 8676 3804 8732
rect 3804 8676 3808 8732
rect 3744 8672 3808 8676
rect 3824 8732 3888 8736
rect 3824 8676 3828 8732
rect 3828 8676 3884 8732
rect 3884 8676 3888 8732
rect 3824 8672 3888 8676
rect 3904 8732 3968 8736
rect 3904 8676 3908 8732
rect 3908 8676 3964 8732
rect 3964 8676 3968 8732
rect 3904 8672 3968 8676
rect 11438 8732 11502 8736
rect 11438 8676 11442 8732
rect 11442 8676 11498 8732
rect 11498 8676 11502 8732
rect 11438 8672 11502 8676
rect 11518 8732 11582 8736
rect 11518 8676 11522 8732
rect 11522 8676 11578 8732
rect 11578 8676 11582 8732
rect 11518 8672 11582 8676
rect 11598 8732 11662 8736
rect 11598 8676 11602 8732
rect 11602 8676 11658 8732
rect 11658 8676 11662 8732
rect 11598 8672 11662 8676
rect 11678 8732 11742 8736
rect 11678 8676 11682 8732
rect 11682 8676 11738 8732
rect 11738 8676 11742 8732
rect 11678 8672 11742 8676
rect 19212 8732 19276 8736
rect 19212 8676 19216 8732
rect 19216 8676 19272 8732
rect 19272 8676 19276 8732
rect 19212 8672 19276 8676
rect 19292 8732 19356 8736
rect 19292 8676 19296 8732
rect 19296 8676 19352 8732
rect 19352 8676 19356 8732
rect 19292 8672 19356 8676
rect 19372 8732 19436 8736
rect 19372 8676 19376 8732
rect 19376 8676 19432 8732
rect 19432 8676 19436 8732
rect 19372 8672 19436 8676
rect 19452 8732 19516 8736
rect 19452 8676 19456 8732
rect 19456 8676 19512 8732
rect 19512 8676 19516 8732
rect 19452 8672 19516 8676
rect 26986 8732 27050 8736
rect 26986 8676 26990 8732
rect 26990 8676 27046 8732
rect 27046 8676 27050 8732
rect 26986 8672 27050 8676
rect 27066 8732 27130 8736
rect 27066 8676 27070 8732
rect 27070 8676 27126 8732
rect 27126 8676 27130 8732
rect 27066 8672 27130 8676
rect 27146 8732 27210 8736
rect 27146 8676 27150 8732
rect 27150 8676 27206 8732
rect 27206 8676 27210 8732
rect 27146 8672 27210 8676
rect 27226 8732 27290 8736
rect 27226 8676 27230 8732
rect 27230 8676 27286 8732
rect 27286 8676 27290 8732
rect 27226 8672 27290 8676
rect 4324 8188 4388 8192
rect 4324 8132 4328 8188
rect 4328 8132 4384 8188
rect 4384 8132 4388 8188
rect 4324 8128 4388 8132
rect 4404 8188 4468 8192
rect 4404 8132 4408 8188
rect 4408 8132 4464 8188
rect 4464 8132 4468 8188
rect 4404 8128 4468 8132
rect 4484 8188 4548 8192
rect 4484 8132 4488 8188
rect 4488 8132 4544 8188
rect 4544 8132 4548 8188
rect 4484 8128 4548 8132
rect 4564 8188 4628 8192
rect 4564 8132 4568 8188
rect 4568 8132 4624 8188
rect 4624 8132 4628 8188
rect 4564 8128 4628 8132
rect 12098 8188 12162 8192
rect 12098 8132 12102 8188
rect 12102 8132 12158 8188
rect 12158 8132 12162 8188
rect 12098 8128 12162 8132
rect 12178 8188 12242 8192
rect 12178 8132 12182 8188
rect 12182 8132 12238 8188
rect 12238 8132 12242 8188
rect 12178 8128 12242 8132
rect 12258 8188 12322 8192
rect 12258 8132 12262 8188
rect 12262 8132 12318 8188
rect 12318 8132 12322 8188
rect 12258 8128 12322 8132
rect 12338 8188 12402 8192
rect 12338 8132 12342 8188
rect 12342 8132 12398 8188
rect 12398 8132 12402 8188
rect 12338 8128 12402 8132
rect 19872 8188 19936 8192
rect 19872 8132 19876 8188
rect 19876 8132 19932 8188
rect 19932 8132 19936 8188
rect 19872 8128 19936 8132
rect 19952 8188 20016 8192
rect 19952 8132 19956 8188
rect 19956 8132 20012 8188
rect 20012 8132 20016 8188
rect 19952 8128 20016 8132
rect 20032 8188 20096 8192
rect 20032 8132 20036 8188
rect 20036 8132 20092 8188
rect 20092 8132 20096 8188
rect 20032 8128 20096 8132
rect 20112 8188 20176 8192
rect 20112 8132 20116 8188
rect 20116 8132 20172 8188
rect 20172 8132 20176 8188
rect 20112 8128 20176 8132
rect 27646 8188 27710 8192
rect 27646 8132 27650 8188
rect 27650 8132 27706 8188
rect 27706 8132 27710 8188
rect 27646 8128 27710 8132
rect 27726 8188 27790 8192
rect 27726 8132 27730 8188
rect 27730 8132 27786 8188
rect 27786 8132 27790 8188
rect 27726 8128 27790 8132
rect 27806 8188 27870 8192
rect 27806 8132 27810 8188
rect 27810 8132 27866 8188
rect 27866 8132 27870 8188
rect 27806 8128 27870 8132
rect 27886 8188 27950 8192
rect 27886 8132 27890 8188
rect 27890 8132 27946 8188
rect 27946 8132 27950 8188
rect 27886 8128 27950 8132
rect 3664 7644 3728 7648
rect 3664 7588 3668 7644
rect 3668 7588 3724 7644
rect 3724 7588 3728 7644
rect 3664 7584 3728 7588
rect 3744 7644 3808 7648
rect 3744 7588 3748 7644
rect 3748 7588 3804 7644
rect 3804 7588 3808 7644
rect 3744 7584 3808 7588
rect 3824 7644 3888 7648
rect 3824 7588 3828 7644
rect 3828 7588 3884 7644
rect 3884 7588 3888 7644
rect 3824 7584 3888 7588
rect 3904 7644 3968 7648
rect 3904 7588 3908 7644
rect 3908 7588 3964 7644
rect 3964 7588 3968 7644
rect 3904 7584 3968 7588
rect 11438 7644 11502 7648
rect 11438 7588 11442 7644
rect 11442 7588 11498 7644
rect 11498 7588 11502 7644
rect 11438 7584 11502 7588
rect 11518 7644 11582 7648
rect 11518 7588 11522 7644
rect 11522 7588 11578 7644
rect 11578 7588 11582 7644
rect 11518 7584 11582 7588
rect 11598 7644 11662 7648
rect 11598 7588 11602 7644
rect 11602 7588 11658 7644
rect 11658 7588 11662 7644
rect 11598 7584 11662 7588
rect 11678 7644 11742 7648
rect 11678 7588 11682 7644
rect 11682 7588 11738 7644
rect 11738 7588 11742 7644
rect 11678 7584 11742 7588
rect 19212 7644 19276 7648
rect 19212 7588 19216 7644
rect 19216 7588 19272 7644
rect 19272 7588 19276 7644
rect 19212 7584 19276 7588
rect 19292 7644 19356 7648
rect 19292 7588 19296 7644
rect 19296 7588 19352 7644
rect 19352 7588 19356 7644
rect 19292 7584 19356 7588
rect 19372 7644 19436 7648
rect 19372 7588 19376 7644
rect 19376 7588 19432 7644
rect 19432 7588 19436 7644
rect 19372 7584 19436 7588
rect 19452 7644 19516 7648
rect 19452 7588 19456 7644
rect 19456 7588 19512 7644
rect 19512 7588 19516 7644
rect 19452 7584 19516 7588
rect 26986 7644 27050 7648
rect 26986 7588 26990 7644
rect 26990 7588 27046 7644
rect 27046 7588 27050 7644
rect 26986 7584 27050 7588
rect 27066 7644 27130 7648
rect 27066 7588 27070 7644
rect 27070 7588 27126 7644
rect 27126 7588 27130 7644
rect 27066 7584 27130 7588
rect 27146 7644 27210 7648
rect 27146 7588 27150 7644
rect 27150 7588 27206 7644
rect 27206 7588 27210 7644
rect 27146 7584 27210 7588
rect 27226 7644 27290 7648
rect 27226 7588 27230 7644
rect 27230 7588 27286 7644
rect 27286 7588 27290 7644
rect 27226 7584 27290 7588
rect 4324 7100 4388 7104
rect 4324 7044 4328 7100
rect 4328 7044 4384 7100
rect 4384 7044 4388 7100
rect 4324 7040 4388 7044
rect 4404 7100 4468 7104
rect 4404 7044 4408 7100
rect 4408 7044 4464 7100
rect 4464 7044 4468 7100
rect 4404 7040 4468 7044
rect 4484 7100 4548 7104
rect 4484 7044 4488 7100
rect 4488 7044 4544 7100
rect 4544 7044 4548 7100
rect 4484 7040 4548 7044
rect 4564 7100 4628 7104
rect 4564 7044 4568 7100
rect 4568 7044 4624 7100
rect 4624 7044 4628 7100
rect 4564 7040 4628 7044
rect 12098 7100 12162 7104
rect 12098 7044 12102 7100
rect 12102 7044 12158 7100
rect 12158 7044 12162 7100
rect 12098 7040 12162 7044
rect 12178 7100 12242 7104
rect 12178 7044 12182 7100
rect 12182 7044 12238 7100
rect 12238 7044 12242 7100
rect 12178 7040 12242 7044
rect 12258 7100 12322 7104
rect 12258 7044 12262 7100
rect 12262 7044 12318 7100
rect 12318 7044 12322 7100
rect 12258 7040 12322 7044
rect 12338 7100 12402 7104
rect 12338 7044 12342 7100
rect 12342 7044 12398 7100
rect 12398 7044 12402 7100
rect 12338 7040 12402 7044
rect 19872 7100 19936 7104
rect 19872 7044 19876 7100
rect 19876 7044 19932 7100
rect 19932 7044 19936 7100
rect 19872 7040 19936 7044
rect 19952 7100 20016 7104
rect 19952 7044 19956 7100
rect 19956 7044 20012 7100
rect 20012 7044 20016 7100
rect 19952 7040 20016 7044
rect 20032 7100 20096 7104
rect 20032 7044 20036 7100
rect 20036 7044 20092 7100
rect 20092 7044 20096 7100
rect 20032 7040 20096 7044
rect 20112 7100 20176 7104
rect 20112 7044 20116 7100
rect 20116 7044 20172 7100
rect 20172 7044 20176 7100
rect 20112 7040 20176 7044
rect 27646 7100 27710 7104
rect 27646 7044 27650 7100
rect 27650 7044 27706 7100
rect 27706 7044 27710 7100
rect 27646 7040 27710 7044
rect 27726 7100 27790 7104
rect 27726 7044 27730 7100
rect 27730 7044 27786 7100
rect 27786 7044 27790 7100
rect 27726 7040 27790 7044
rect 27806 7100 27870 7104
rect 27806 7044 27810 7100
rect 27810 7044 27866 7100
rect 27866 7044 27870 7100
rect 27806 7040 27870 7044
rect 27886 7100 27950 7104
rect 27886 7044 27890 7100
rect 27890 7044 27946 7100
rect 27946 7044 27950 7100
rect 27886 7040 27950 7044
rect 3664 6556 3728 6560
rect 3664 6500 3668 6556
rect 3668 6500 3724 6556
rect 3724 6500 3728 6556
rect 3664 6496 3728 6500
rect 3744 6556 3808 6560
rect 3744 6500 3748 6556
rect 3748 6500 3804 6556
rect 3804 6500 3808 6556
rect 3744 6496 3808 6500
rect 3824 6556 3888 6560
rect 3824 6500 3828 6556
rect 3828 6500 3884 6556
rect 3884 6500 3888 6556
rect 3824 6496 3888 6500
rect 3904 6556 3968 6560
rect 3904 6500 3908 6556
rect 3908 6500 3964 6556
rect 3964 6500 3968 6556
rect 3904 6496 3968 6500
rect 11438 6556 11502 6560
rect 11438 6500 11442 6556
rect 11442 6500 11498 6556
rect 11498 6500 11502 6556
rect 11438 6496 11502 6500
rect 11518 6556 11582 6560
rect 11518 6500 11522 6556
rect 11522 6500 11578 6556
rect 11578 6500 11582 6556
rect 11518 6496 11582 6500
rect 11598 6556 11662 6560
rect 11598 6500 11602 6556
rect 11602 6500 11658 6556
rect 11658 6500 11662 6556
rect 11598 6496 11662 6500
rect 11678 6556 11742 6560
rect 11678 6500 11682 6556
rect 11682 6500 11738 6556
rect 11738 6500 11742 6556
rect 11678 6496 11742 6500
rect 19212 6556 19276 6560
rect 19212 6500 19216 6556
rect 19216 6500 19272 6556
rect 19272 6500 19276 6556
rect 19212 6496 19276 6500
rect 19292 6556 19356 6560
rect 19292 6500 19296 6556
rect 19296 6500 19352 6556
rect 19352 6500 19356 6556
rect 19292 6496 19356 6500
rect 19372 6556 19436 6560
rect 19372 6500 19376 6556
rect 19376 6500 19432 6556
rect 19432 6500 19436 6556
rect 19372 6496 19436 6500
rect 19452 6556 19516 6560
rect 19452 6500 19456 6556
rect 19456 6500 19512 6556
rect 19512 6500 19516 6556
rect 19452 6496 19516 6500
rect 26986 6556 27050 6560
rect 26986 6500 26990 6556
rect 26990 6500 27046 6556
rect 27046 6500 27050 6556
rect 26986 6496 27050 6500
rect 27066 6556 27130 6560
rect 27066 6500 27070 6556
rect 27070 6500 27126 6556
rect 27126 6500 27130 6556
rect 27066 6496 27130 6500
rect 27146 6556 27210 6560
rect 27146 6500 27150 6556
rect 27150 6500 27206 6556
rect 27206 6500 27210 6556
rect 27146 6496 27210 6500
rect 27226 6556 27290 6560
rect 27226 6500 27230 6556
rect 27230 6500 27286 6556
rect 27286 6500 27290 6556
rect 27226 6496 27290 6500
rect 4324 6012 4388 6016
rect 4324 5956 4328 6012
rect 4328 5956 4384 6012
rect 4384 5956 4388 6012
rect 4324 5952 4388 5956
rect 4404 6012 4468 6016
rect 4404 5956 4408 6012
rect 4408 5956 4464 6012
rect 4464 5956 4468 6012
rect 4404 5952 4468 5956
rect 4484 6012 4548 6016
rect 4484 5956 4488 6012
rect 4488 5956 4544 6012
rect 4544 5956 4548 6012
rect 4484 5952 4548 5956
rect 4564 6012 4628 6016
rect 4564 5956 4568 6012
rect 4568 5956 4624 6012
rect 4624 5956 4628 6012
rect 4564 5952 4628 5956
rect 12098 6012 12162 6016
rect 12098 5956 12102 6012
rect 12102 5956 12158 6012
rect 12158 5956 12162 6012
rect 12098 5952 12162 5956
rect 12178 6012 12242 6016
rect 12178 5956 12182 6012
rect 12182 5956 12238 6012
rect 12238 5956 12242 6012
rect 12178 5952 12242 5956
rect 12258 6012 12322 6016
rect 12258 5956 12262 6012
rect 12262 5956 12318 6012
rect 12318 5956 12322 6012
rect 12258 5952 12322 5956
rect 12338 6012 12402 6016
rect 12338 5956 12342 6012
rect 12342 5956 12398 6012
rect 12398 5956 12402 6012
rect 12338 5952 12402 5956
rect 19872 6012 19936 6016
rect 19872 5956 19876 6012
rect 19876 5956 19932 6012
rect 19932 5956 19936 6012
rect 19872 5952 19936 5956
rect 19952 6012 20016 6016
rect 19952 5956 19956 6012
rect 19956 5956 20012 6012
rect 20012 5956 20016 6012
rect 19952 5952 20016 5956
rect 20032 6012 20096 6016
rect 20032 5956 20036 6012
rect 20036 5956 20092 6012
rect 20092 5956 20096 6012
rect 20032 5952 20096 5956
rect 20112 6012 20176 6016
rect 20112 5956 20116 6012
rect 20116 5956 20172 6012
rect 20172 5956 20176 6012
rect 20112 5952 20176 5956
rect 27646 6012 27710 6016
rect 27646 5956 27650 6012
rect 27650 5956 27706 6012
rect 27706 5956 27710 6012
rect 27646 5952 27710 5956
rect 27726 6012 27790 6016
rect 27726 5956 27730 6012
rect 27730 5956 27786 6012
rect 27786 5956 27790 6012
rect 27726 5952 27790 5956
rect 27806 6012 27870 6016
rect 27806 5956 27810 6012
rect 27810 5956 27866 6012
rect 27866 5956 27870 6012
rect 27806 5952 27870 5956
rect 27886 6012 27950 6016
rect 27886 5956 27890 6012
rect 27890 5956 27946 6012
rect 27946 5956 27950 6012
rect 27886 5952 27950 5956
rect 3664 5468 3728 5472
rect 3664 5412 3668 5468
rect 3668 5412 3724 5468
rect 3724 5412 3728 5468
rect 3664 5408 3728 5412
rect 3744 5468 3808 5472
rect 3744 5412 3748 5468
rect 3748 5412 3804 5468
rect 3804 5412 3808 5468
rect 3744 5408 3808 5412
rect 3824 5468 3888 5472
rect 3824 5412 3828 5468
rect 3828 5412 3884 5468
rect 3884 5412 3888 5468
rect 3824 5408 3888 5412
rect 3904 5468 3968 5472
rect 3904 5412 3908 5468
rect 3908 5412 3964 5468
rect 3964 5412 3968 5468
rect 3904 5408 3968 5412
rect 11438 5468 11502 5472
rect 11438 5412 11442 5468
rect 11442 5412 11498 5468
rect 11498 5412 11502 5468
rect 11438 5408 11502 5412
rect 11518 5468 11582 5472
rect 11518 5412 11522 5468
rect 11522 5412 11578 5468
rect 11578 5412 11582 5468
rect 11518 5408 11582 5412
rect 11598 5468 11662 5472
rect 11598 5412 11602 5468
rect 11602 5412 11658 5468
rect 11658 5412 11662 5468
rect 11598 5408 11662 5412
rect 11678 5468 11742 5472
rect 11678 5412 11682 5468
rect 11682 5412 11738 5468
rect 11738 5412 11742 5468
rect 11678 5408 11742 5412
rect 19212 5468 19276 5472
rect 19212 5412 19216 5468
rect 19216 5412 19272 5468
rect 19272 5412 19276 5468
rect 19212 5408 19276 5412
rect 19292 5468 19356 5472
rect 19292 5412 19296 5468
rect 19296 5412 19352 5468
rect 19352 5412 19356 5468
rect 19292 5408 19356 5412
rect 19372 5468 19436 5472
rect 19372 5412 19376 5468
rect 19376 5412 19432 5468
rect 19432 5412 19436 5468
rect 19372 5408 19436 5412
rect 19452 5468 19516 5472
rect 19452 5412 19456 5468
rect 19456 5412 19512 5468
rect 19512 5412 19516 5468
rect 19452 5408 19516 5412
rect 26986 5468 27050 5472
rect 26986 5412 26990 5468
rect 26990 5412 27046 5468
rect 27046 5412 27050 5468
rect 26986 5408 27050 5412
rect 27066 5468 27130 5472
rect 27066 5412 27070 5468
rect 27070 5412 27126 5468
rect 27126 5412 27130 5468
rect 27066 5408 27130 5412
rect 27146 5468 27210 5472
rect 27146 5412 27150 5468
rect 27150 5412 27206 5468
rect 27206 5412 27210 5468
rect 27146 5408 27210 5412
rect 27226 5468 27290 5472
rect 27226 5412 27230 5468
rect 27230 5412 27286 5468
rect 27286 5412 27290 5468
rect 27226 5408 27290 5412
rect 4324 4924 4388 4928
rect 4324 4868 4328 4924
rect 4328 4868 4384 4924
rect 4384 4868 4388 4924
rect 4324 4864 4388 4868
rect 4404 4924 4468 4928
rect 4404 4868 4408 4924
rect 4408 4868 4464 4924
rect 4464 4868 4468 4924
rect 4404 4864 4468 4868
rect 4484 4924 4548 4928
rect 4484 4868 4488 4924
rect 4488 4868 4544 4924
rect 4544 4868 4548 4924
rect 4484 4864 4548 4868
rect 4564 4924 4628 4928
rect 4564 4868 4568 4924
rect 4568 4868 4624 4924
rect 4624 4868 4628 4924
rect 4564 4864 4628 4868
rect 12098 4924 12162 4928
rect 12098 4868 12102 4924
rect 12102 4868 12158 4924
rect 12158 4868 12162 4924
rect 12098 4864 12162 4868
rect 12178 4924 12242 4928
rect 12178 4868 12182 4924
rect 12182 4868 12238 4924
rect 12238 4868 12242 4924
rect 12178 4864 12242 4868
rect 12258 4924 12322 4928
rect 12258 4868 12262 4924
rect 12262 4868 12318 4924
rect 12318 4868 12322 4924
rect 12258 4864 12322 4868
rect 12338 4924 12402 4928
rect 12338 4868 12342 4924
rect 12342 4868 12398 4924
rect 12398 4868 12402 4924
rect 12338 4864 12402 4868
rect 19872 4924 19936 4928
rect 19872 4868 19876 4924
rect 19876 4868 19932 4924
rect 19932 4868 19936 4924
rect 19872 4864 19936 4868
rect 19952 4924 20016 4928
rect 19952 4868 19956 4924
rect 19956 4868 20012 4924
rect 20012 4868 20016 4924
rect 19952 4864 20016 4868
rect 20032 4924 20096 4928
rect 20032 4868 20036 4924
rect 20036 4868 20092 4924
rect 20092 4868 20096 4924
rect 20032 4864 20096 4868
rect 20112 4924 20176 4928
rect 20112 4868 20116 4924
rect 20116 4868 20172 4924
rect 20172 4868 20176 4924
rect 20112 4864 20176 4868
rect 27646 4924 27710 4928
rect 27646 4868 27650 4924
rect 27650 4868 27706 4924
rect 27706 4868 27710 4924
rect 27646 4864 27710 4868
rect 27726 4924 27790 4928
rect 27726 4868 27730 4924
rect 27730 4868 27786 4924
rect 27786 4868 27790 4924
rect 27726 4864 27790 4868
rect 27806 4924 27870 4928
rect 27806 4868 27810 4924
rect 27810 4868 27866 4924
rect 27866 4868 27870 4924
rect 27806 4864 27870 4868
rect 27886 4924 27950 4928
rect 27886 4868 27890 4924
rect 27890 4868 27946 4924
rect 27946 4868 27950 4924
rect 27886 4864 27950 4868
rect 3664 4380 3728 4384
rect 3664 4324 3668 4380
rect 3668 4324 3724 4380
rect 3724 4324 3728 4380
rect 3664 4320 3728 4324
rect 3744 4380 3808 4384
rect 3744 4324 3748 4380
rect 3748 4324 3804 4380
rect 3804 4324 3808 4380
rect 3744 4320 3808 4324
rect 3824 4380 3888 4384
rect 3824 4324 3828 4380
rect 3828 4324 3884 4380
rect 3884 4324 3888 4380
rect 3824 4320 3888 4324
rect 3904 4380 3968 4384
rect 3904 4324 3908 4380
rect 3908 4324 3964 4380
rect 3964 4324 3968 4380
rect 3904 4320 3968 4324
rect 11438 4380 11502 4384
rect 11438 4324 11442 4380
rect 11442 4324 11498 4380
rect 11498 4324 11502 4380
rect 11438 4320 11502 4324
rect 11518 4380 11582 4384
rect 11518 4324 11522 4380
rect 11522 4324 11578 4380
rect 11578 4324 11582 4380
rect 11518 4320 11582 4324
rect 11598 4380 11662 4384
rect 11598 4324 11602 4380
rect 11602 4324 11658 4380
rect 11658 4324 11662 4380
rect 11598 4320 11662 4324
rect 11678 4380 11742 4384
rect 11678 4324 11682 4380
rect 11682 4324 11738 4380
rect 11738 4324 11742 4380
rect 11678 4320 11742 4324
rect 19212 4380 19276 4384
rect 19212 4324 19216 4380
rect 19216 4324 19272 4380
rect 19272 4324 19276 4380
rect 19212 4320 19276 4324
rect 19292 4380 19356 4384
rect 19292 4324 19296 4380
rect 19296 4324 19352 4380
rect 19352 4324 19356 4380
rect 19292 4320 19356 4324
rect 19372 4380 19436 4384
rect 19372 4324 19376 4380
rect 19376 4324 19432 4380
rect 19432 4324 19436 4380
rect 19372 4320 19436 4324
rect 19452 4380 19516 4384
rect 19452 4324 19456 4380
rect 19456 4324 19512 4380
rect 19512 4324 19516 4380
rect 19452 4320 19516 4324
rect 26986 4380 27050 4384
rect 26986 4324 26990 4380
rect 26990 4324 27046 4380
rect 27046 4324 27050 4380
rect 26986 4320 27050 4324
rect 27066 4380 27130 4384
rect 27066 4324 27070 4380
rect 27070 4324 27126 4380
rect 27126 4324 27130 4380
rect 27066 4320 27130 4324
rect 27146 4380 27210 4384
rect 27146 4324 27150 4380
rect 27150 4324 27206 4380
rect 27206 4324 27210 4380
rect 27146 4320 27210 4324
rect 27226 4380 27290 4384
rect 27226 4324 27230 4380
rect 27230 4324 27286 4380
rect 27286 4324 27290 4380
rect 27226 4320 27290 4324
rect 4324 3836 4388 3840
rect 4324 3780 4328 3836
rect 4328 3780 4384 3836
rect 4384 3780 4388 3836
rect 4324 3776 4388 3780
rect 4404 3836 4468 3840
rect 4404 3780 4408 3836
rect 4408 3780 4464 3836
rect 4464 3780 4468 3836
rect 4404 3776 4468 3780
rect 4484 3836 4548 3840
rect 4484 3780 4488 3836
rect 4488 3780 4544 3836
rect 4544 3780 4548 3836
rect 4484 3776 4548 3780
rect 4564 3836 4628 3840
rect 4564 3780 4568 3836
rect 4568 3780 4624 3836
rect 4624 3780 4628 3836
rect 4564 3776 4628 3780
rect 12098 3836 12162 3840
rect 12098 3780 12102 3836
rect 12102 3780 12158 3836
rect 12158 3780 12162 3836
rect 12098 3776 12162 3780
rect 12178 3836 12242 3840
rect 12178 3780 12182 3836
rect 12182 3780 12238 3836
rect 12238 3780 12242 3836
rect 12178 3776 12242 3780
rect 12258 3836 12322 3840
rect 12258 3780 12262 3836
rect 12262 3780 12318 3836
rect 12318 3780 12322 3836
rect 12258 3776 12322 3780
rect 12338 3836 12402 3840
rect 12338 3780 12342 3836
rect 12342 3780 12398 3836
rect 12398 3780 12402 3836
rect 12338 3776 12402 3780
rect 19872 3836 19936 3840
rect 19872 3780 19876 3836
rect 19876 3780 19932 3836
rect 19932 3780 19936 3836
rect 19872 3776 19936 3780
rect 19952 3836 20016 3840
rect 19952 3780 19956 3836
rect 19956 3780 20012 3836
rect 20012 3780 20016 3836
rect 19952 3776 20016 3780
rect 20032 3836 20096 3840
rect 20032 3780 20036 3836
rect 20036 3780 20092 3836
rect 20092 3780 20096 3836
rect 20032 3776 20096 3780
rect 20112 3836 20176 3840
rect 20112 3780 20116 3836
rect 20116 3780 20172 3836
rect 20172 3780 20176 3836
rect 20112 3776 20176 3780
rect 27646 3836 27710 3840
rect 27646 3780 27650 3836
rect 27650 3780 27706 3836
rect 27706 3780 27710 3836
rect 27646 3776 27710 3780
rect 27726 3836 27790 3840
rect 27726 3780 27730 3836
rect 27730 3780 27786 3836
rect 27786 3780 27790 3836
rect 27726 3776 27790 3780
rect 27806 3836 27870 3840
rect 27806 3780 27810 3836
rect 27810 3780 27866 3836
rect 27866 3780 27870 3836
rect 27806 3776 27870 3780
rect 27886 3836 27950 3840
rect 27886 3780 27890 3836
rect 27890 3780 27946 3836
rect 27946 3780 27950 3836
rect 27886 3776 27950 3780
rect 3664 3292 3728 3296
rect 3664 3236 3668 3292
rect 3668 3236 3724 3292
rect 3724 3236 3728 3292
rect 3664 3232 3728 3236
rect 3744 3292 3808 3296
rect 3744 3236 3748 3292
rect 3748 3236 3804 3292
rect 3804 3236 3808 3292
rect 3744 3232 3808 3236
rect 3824 3292 3888 3296
rect 3824 3236 3828 3292
rect 3828 3236 3884 3292
rect 3884 3236 3888 3292
rect 3824 3232 3888 3236
rect 3904 3292 3968 3296
rect 3904 3236 3908 3292
rect 3908 3236 3964 3292
rect 3964 3236 3968 3292
rect 3904 3232 3968 3236
rect 11438 3292 11502 3296
rect 11438 3236 11442 3292
rect 11442 3236 11498 3292
rect 11498 3236 11502 3292
rect 11438 3232 11502 3236
rect 11518 3292 11582 3296
rect 11518 3236 11522 3292
rect 11522 3236 11578 3292
rect 11578 3236 11582 3292
rect 11518 3232 11582 3236
rect 11598 3292 11662 3296
rect 11598 3236 11602 3292
rect 11602 3236 11658 3292
rect 11658 3236 11662 3292
rect 11598 3232 11662 3236
rect 11678 3292 11742 3296
rect 11678 3236 11682 3292
rect 11682 3236 11738 3292
rect 11738 3236 11742 3292
rect 11678 3232 11742 3236
rect 19212 3292 19276 3296
rect 19212 3236 19216 3292
rect 19216 3236 19272 3292
rect 19272 3236 19276 3292
rect 19212 3232 19276 3236
rect 19292 3292 19356 3296
rect 19292 3236 19296 3292
rect 19296 3236 19352 3292
rect 19352 3236 19356 3292
rect 19292 3232 19356 3236
rect 19372 3292 19436 3296
rect 19372 3236 19376 3292
rect 19376 3236 19432 3292
rect 19432 3236 19436 3292
rect 19372 3232 19436 3236
rect 19452 3292 19516 3296
rect 19452 3236 19456 3292
rect 19456 3236 19512 3292
rect 19512 3236 19516 3292
rect 19452 3232 19516 3236
rect 26986 3292 27050 3296
rect 26986 3236 26990 3292
rect 26990 3236 27046 3292
rect 27046 3236 27050 3292
rect 26986 3232 27050 3236
rect 27066 3292 27130 3296
rect 27066 3236 27070 3292
rect 27070 3236 27126 3292
rect 27126 3236 27130 3292
rect 27066 3232 27130 3236
rect 27146 3292 27210 3296
rect 27146 3236 27150 3292
rect 27150 3236 27206 3292
rect 27206 3236 27210 3292
rect 27146 3232 27210 3236
rect 27226 3292 27290 3296
rect 27226 3236 27230 3292
rect 27230 3236 27286 3292
rect 27286 3236 27290 3292
rect 27226 3232 27290 3236
rect 4324 2748 4388 2752
rect 4324 2692 4328 2748
rect 4328 2692 4384 2748
rect 4384 2692 4388 2748
rect 4324 2688 4388 2692
rect 4404 2748 4468 2752
rect 4404 2692 4408 2748
rect 4408 2692 4464 2748
rect 4464 2692 4468 2748
rect 4404 2688 4468 2692
rect 4484 2748 4548 2752
rect 4484 2692 4488 2748
rect 4488 2692 4544 2748
rect 4544 2692 4548 2748
rect 4484 2688 4548 2692
rect 4564 2748 4628 2752
rect 4564 2692 4568 2748
rect 4568 2692 4624 2748
rect 4624 2692 4628 2748
rect 4564 2688 4628 2692
rect 12098 2748 12162 2752
rect 12098 2692 12102 2748
rect 12102 2692 12158 2748
rect 12158 2692 12162 2748
rect 12098 2688 12162 2692
rect 12178 2748 12242 2752
rect 12178 2692 12182 2748
rect 12182 2692 12238 2748
rect 12238 2692 12242 2748
rect 12178 2688 12242 2692
rect 12258 2748 12322 2752
rect 12258 2692 12262 2748
rect 12262 2692 12318 2748
rect 12318 2692 12322 2748
rect 12258 2688 12322 2692
rect 12338 2748 12402 2752
rect 12338 2692 12342 2748
rect 12342 2692 12398 2748
rect 12398 2692 12402 2748
rect 12338 2688 12402 2692
rect 19872 2748 19936 2752
rect 19872 2692 19876 2748
rect 19876 2692 19932 2748
rect 19932 2692 19936 2748
rect 19872 2688 19936 2692
rect 19952 2748 20016 2752
rect 19952 2692 19956 2748
rect 19956 2692 20012 2748
rect 20012 2692 20016 2748
rect 19952 2688 20016 2692
rect 20032 2748 20096 2752
rect 20032 2692 20036 2748
rect 20036 2692 20092 2748
rect 20092 2692 20096 2748
rect 20032 2688 20096 2692
rect 20112 2748 20176 2752
rect 20112 2692 20116 2748
rect 20116 2692 20172 2748
rect 20172 2692 20176 2748
rect 20112 2688 20176 2692
rect 27646 2748 27710 2752
rect 27646 2692 27650 2748
rect 27650 2692 27706 2748
rect 27706 2692 27710 2748
rect 27646 2688 27710 2692
rect 27726 2748 27790 2752
rect 27726 2692 27730 2748
rect 27730 2692 27786 2748
rect 27786 2692 27790 2748
rect 27726 2688 27790 2692
rect 27806 2748 27870 2752
rect 27806 2692 27810 2748
rect 27810 2692 27866 2748
rect 27866 2692 27870 2748
rect 27806 2688 27870 2692
rect 27886 2748 27950 2752
rect 27886 2692 27890 2748
rect 27890 2692 27946 2748
rect 27946 2692 27950 2748
rect 27886 2688 27950 2692
rect 3664 2204 3728 2208
rect 3664 2148 3668 2204
rect 3668 2148 3724 2204
rect 3724 2148 3728 2204
rect 3664 2144 3728 2148
rect 3744 2204 3808 2208
rect 3744 2148 3748 2204
rect 3748 2148 3804 2204
rect 3804 2148 3808 2204
rect 3744 2144 3808 2148
rect 3824 2204 3888 2208
rect 3824 2148 3828 2204
rect 3828 2148 3884 2204
rect 3884 2148 3888 2204
rect 3824 2144 3888 2148
rect 3904 2204 3968 2208
rect 3904 2148 3908 2204
rect 3908 2148 3964 2204
rect 3964 2148 3968 2204
rect 3904 2144 3968 2148
rect 11438 2204 11502 2208
rect 11438 2148 11442 2204
rect 11442 2148 11498 2204
rect 11498 2148 11502 2204
rect 11438 2144 11502 2148
rect 11518 2204 11582 2208
rect 11518 2148 11522 2204
rect 11522 2148 11578 2204
rect 11578 2148 11582 2204
rect 11518 2144 11582 2148
rect 11598 2204 11662 2208
rect 11598 2148 11602 2204
rect 11602 2148 11658 2204
rect 11658 2148 11662 2204
rect 11598 2144 11662 2148
rect 11678 2204 11742 2208
rect 11678 2148 11682 2204
rect 11682 2148 11738 2204
rect 11738 2148 11742 2204
rect 11678 2144 11742 2148
rect 19212 2204 19276 2208
rect 19212 2148 19216 2204
rect 19216 2148 19272 2204
rect 19272 2148 19276 2204
rect 19212 2144 19276 2148
rect 19292 2204 19356 2208
rect 19292 2148 19296 2204
rect 19296 2148 19352 2204
rect 19352 2148 19356 2204
rect 19292 2144 19356 2148
rect 19372 2204 19436 2208
rect 19372 2148 19376 2204
rect 19376 2148 19432 2204
rect 19432 2148 19436 2204
rect 19372 2144 19436 2148
rect 19452 2204 19516 2208
rect 19452 2148 19456 2204
rect 19456 2148 19512 2204
rect 19512 2148 19516 2204
rect 19452 2144 19516 2148
rect 26986 2204 27050 2208
rect 26986 2148 26990 2204
rect 26990 2148 27046 2204
rect 27046 2148 27050 2204
rect 26986 2144 27050 2148
rect 27066 2204 27130 2208
rect 27066 2148 27070 2204
rect 27070 2148 27126 2204
rect 27126 2148 27130 2204
rect 27066 2144 27130 2148
rect 27146 2204 27210 2208
rect 27146 2148 27150 2204
rect 27150 2148 27206 2204
rect 27206 2148 27210 2204
rect 27146 2144 27210 2148
rect 27226 2204 27290 2208
rect 27226 2148 27230 2204
rect 27230 2148 27286 2204
rect 27286 2148 27290 2204
rect 27226 2144 27290 2148
rect 4324 1660 4388 1664
rect 4324 1604 4328 1660
rect 4328 1604 4384 1660
rect 4384 1604 4388 1660
rect 4324 1600 4388 1604
rect 4404 1660 4468 1664
rect 4404 1604 4408 1660
rect 4408 1604 4464 1660
rect 4464 1604 4468 1660
rect 4404 1600 4468 1604
rect 4484 1660 4548 1664
rect 4484 1604 4488 1660
rect 4488 1604 4544 1660
rect 4544 1604 4548 1660
rect 4484 1600 4548 1604
rect 4564 1660 4628 1664
rect 4564 1604 4568 1660
rect 4568 1604 4624 1660
rect 4624 1604 4628 1660
rect 4564 1600 4628 1604
rect 12098 1660 12162 1664
rect 12098 1604 12102 1660
rect 12102 1604 12158 1660
rect 12158 1604 12162 1660
rect 12098 1600 12162 1604
rect 12178 1660 12242 1664
rect 12178 1604 12182 1660
rect 12182 1604 12238 1660
rect 12238 1604 12242 1660
rect 12178 1600 12242 1604
rect 12258 1660 12322 1664
rect 12258 1604 12262 1660
rect 12262 1604 12318 1660
rect 12318 1604 12322 1660
rect 12258 1600 12322 1604
rect 12338 1660 12402 1664
rect 12338 1604 12342 1660
rect 12342 1604 12398 1660
rect 12398 1604 12402 1660
rect 12338 1600 12402 1604
rect 19872 1660 19936 1664
rect 19872 1604 19876 1660
rect 19876 1604 19932 1660
rect 19932 1604 19936 1660
rect 19872 1600 19936 1604
rect 19952 1660 20016 1664
rect 19952 1604 19956 1660
rect 19956 1604 20012 1660
rect 20012 1604 20016 1660
rect 19952 1600 20016 1604
rect 20032 1660 20096 1664
rect 20032 1604 20036 1660
rect 20036 1604 20092 1660
rect 20092 1604 20096 1660
rect 20032 1600 20096 1604
rect 20112 1660 20176 1664
rect 20112 1604 20116 1660
rect 20116 1604 20172 1660
rect 20172 1604 20176 1660
rect 20112 1600 20176 1604
rect 27646 1660 27710 1664
rect 27646 1604 27650 1660
rect 27650 1604 27706 1660
rect 27706 1604 27710 1660
rect 27646 1600 27710 1604
rect 27726 1660 27790 1664
rect 27726 1604 27730 1660
rect 27730 1604 27786 1660
rect 27786 1604 27790 1660
rect 27726 1600 27790 1604
rect 27806 1660 27870 1664
rect 27806 1604 27810 1660
rect 27810 1604 27866 1660
rect 27866 1604 27870 1660
rect 27806 1600 27870 1604
rect 27886 1660 27950 1664
rect 27886 1604 27890 1660
rect 27890 1604 27946 1660
rect 27946 1604 27950 1660
rect 27886 1600 27950 1604
rect 3664 1116 3728 1120
rect 3664 1060 3668 1116
rect 3668 1060 3724 1116
rect 3724 1060 3728 1116
rect 3664 1056 3728 1060
rect 3744 1116 3808 1120
rect 3744 1060 3748 1116
rect 3748 1060 3804 1116
rect 3804 1060 3808 1116
rect 3744 1056 3808 1060
rect 3824 1116 3888 1120
rect 3824 1060 3828 1116
rect 3828 1060 3884 1116
rect 3884 1060 3888 1116
rect 3824 1056 3888 1060
rect 3904 1116 3968 1120
rect 3904 1060 3908 1116
rect 3908 1060 3964 1116
rect 3964 1060 3968 1116
rect 3904 1056 3968 1060
rect 11438 1116 11502 1120
rect 11438 1060 11442 1116
rect 11442 1060 11498 1116
rect 11498 1060 11502 1116
rect 11438 1056 11502 1060
rect 11518 1116 11582 1120
rect 11518 1060 11522 1116
rect 11522 1060 11578 1116
rect 11578 1060 11582 1116
rect 11518 1056 11582 1060
rect 11598 1116 11662 1120
rect 11598 1060 11602 1116
rect 11602 1060 11658 1116
rect 11658 1060 11662 1116
rect 11598 1056 11662 1060
rect 11678 1116 11742 1120
rect 11678 1060 11682 1116
rect 11682 1060 11738 1116
rect 11738 1060 11742 1116
rect 11678 1056 11742 1060
rect 19212 1116 19276 1120
rect 19212 1060 19216 1116
rect 19216 1060 19272 1116
rect 19272 1060 19276 1116
rect 19212 1056 19276 1060
rect 19292 1116 19356 1120
rect 19292 1060 19296 1116
rect 19296 1060 19352 1116
rect 19352 1060 19356 1116
rect 19292 1056 19356 1060
rect 19372 1116 19436 1120
rect 19372 1060 19376 1116
rect 19376 1060 19432 1116
rect 19432 1060 19436 1116
rect 19372 1056 19436 1060
rect 19452 1116 19516 1120
rect 19452 1060 19456 1116
rect 19456 1060 19512 1116
rect 19512 1060 19516 1116
rect 19452 1056 19516 1060
rect 26986 1116 27050 1120
rect 26986 1060 26990 1116
rect 26990 1060 27046 1116
rect 27046 1060 27050 1116
rect 26986 1056 27050 1060
rect 27066 1116 27130 1120
rect 27066 1060 27070 1116
rect 27070 1060 27126 1116
rect 27126 1060 27130 1116
rect 27066 1056 27130 1060
rect 27146 1116 27210 1120
rect 27146 1060 27150 1116
rect 27150 1060 27206 1116
rect 27206 1060 27210 1116
rect 27146 1056 27210 1060
rect 27226 1116 27290 1120
rect 27226 1060 27230 1116
rect 27230 1060 27286 1116
rect 27286 1060 27290 1116
rect 27226 1056 27290 1060
rect 4324 572 4388 576
rect 4324 516 4328 572
rect 4328 516 4384 572
rect 4384 516 4388 572
rect 4324 512 4388 516
rect 4404 572 4468 576
rect 4404 516 4408 572
rect 4408 516 4464 572
rect 4464 516 4468 572
rect 4404 512 4468 516
rect 4484 572 4548 576
rect 4484 516 4488 572
rect 4488 516 4544 572
rect 4544 516 4548 572
rect 4484 512 4548 516
rect 4564 572 4628 576
rect 4564 516 4568 572
rect 4568 516 4624 572
rect 4624 516 4628 572
rect 4564 512 4628 516
rect 12098 572 12162 576
rect 12098 516 12102 572
rect 12102 516 12158 572
rect 12158 516 12162 572
rect 12098 512 12162 516
rect 12178 572 12242 576
rect 12178 516 12182 572
rect 12182 516 12238 572
rect 12238 516 12242 572
rect 12178 512 12242 516
rect 12258 572 12322 576
rect 12258 516 12262 572
rect 12262 516 12318 572
rect 12318 516 12322 572
rect 12258 512 12322 516
rect 12338 572 12402 576
rect 12338 516 12342 572
rect 12342 516 12398 572
rect 12398 516 12402 572
rect 12338 512 12402 516
rect 19872 572 19936 576
rect 19872 516 19876 572
rect 19876 516 19932 572
rect 19932 516 19936 572
rect 19872 512 19936 516
rect 19952 572 20016 576
rect 19952 516 19956 572
rect 19956 516 20012 572
rect 20012 516 20016 572
rect 19952 512 20016 516
rect 20032 572 20096 576
rect 20032 516 20036 572
rect 20036 516 20092 572
rect 20092 516 20096 572
rect 20032 512 20096 516
rect 20112 572 20176 576
rect 20112 516 20116 572
rect 20116 516 20172 572
rect 20172 516 20176 572
rect 20112 512 20176 516
rect 27646 572 27710 576
rect 27646 516 27650 572
rect 27650 516 27706 572
rect 27706 516 27710 572
rect 27646 512 27710 516
rect 27726 572 27790 576
rect 27726 516 27730 572
rect 27730 516 27786 572
rect 27786 516 27790 572
rect 27726 512 27790 516
rect 27806 572 27870 576
rect 27806 516 27810 572
rect 27810 516 27866 572
rect 27866 516 27870 572
rect 27806 512 27870 516
rect 27886 572 27950 576
rect 27886 516 27890 572
rect 27890 516 27946 572
rect 27946 516 27950 572
rect 27886 512 27950 516
<< metal4 >>
rect 3656 18528 3976 19088
rect 3656 18464 3664 18528
rect 3728 18464 3744 18528
rect 3808 18464 3824 18528
rect 3888 18464 3904 18528
rect 3968 18464 3976 18528
rect 3656 17440 3976 18464
rect 3656 17376 3664 17440
rect 3728 17376 3744 17440
rect 3808 17376 3824 17440
rect 3888 17376 3904 17440
rect 3968 17376 3976 17440
rect 3656 16352 3976 17376
rect 3656 16288 3664 16352
rect 3728 16288 3744 16352
rect 3808 16288 3824 16352
rect 3888 16288 3904 16352
rect 3968 16288 3976 16352
rect 3656 15264 3976 16288
rect 3656 15200 3664 15264
rect 3728 15200 3744 15264
rect 3808 15200 3824 15264
rect 3888 15200 3904 15264
rect 3968 15200 3976 15264
rect 3656 14176 3976 15200
rect 3656 14112 3664 14176
rect 3728 14112 3744 14176
rect 3808 14112 3824 14176
rect 3888 14112 3904 14176
rect 3968 14112 3976 14176
rect 3656 13088 3976 14112
rect 3656 13024 3664 13088
rect 3728 13024 3744 13088
rect 3808 13024 3824 13088
rect 3888 13024 3904 13088
rect 3968 13024 3976 13088
rect 3656 12000 3976 13024
rect 3656 11936 3664 12000
rect 3728 11936 3744 12000
rect 3808 11936 3824 12000
rect 3888 11936 3904 12000
rect 3968 11936 3976 12000
rect 3656 10912 3976 11936
rect 3656 10848 3664 10912
rect 3728 10848 3744 10912
rect 3808 10848 3824 10912
rect 3888 10848 3904 10912
rect 3968 10848 3976 10912
rect 3656 9824 3976 10848
rect 3656 9760 3664 9824
rect 3728 9760 3744 9824
rect 3808 9760 3824 9824
rect 3888 9760 3904 9824
rect 3968 9760 3976 9824
rect 3656 8736 3976 9760
rect 3656 8672 3664 8736
rect 3728 8672 3744 8736
rect 3808 8672 3824 8736
rect 3888 8672 3904 8736
rect 3968 8672 3976 8736
rect 3656 7648 3976 8672
rect 3656 7584 3664 7648
rect 3728 7584 3744 7648
rect 3808 7584 3824 7648
rect 3888 7584 3904 7648
rect 3968 7584 3976 7648
rect 3656 6560 3976 7584
rect 3656 6496 3664 6560
rect 3728 6496 3744 6560
rect 3808 6496 3824 6560
rect 3888 6496 3904 6560
rect 3968 6496 3976 6560
rect 3656 5472 3976 6496
rect 3656 5408 3664 5472
rect 3728 5408 3744 5472
rect 3808 5408 3824 5472
rect 3888 5408 3904 5472
rect 3968 5408 3976 5472
rect 3656 4384 3976 5408
rect 3656 4320 3664 4384
rect 3728 4320 3744 4384
rect 3808 4320 3824 4384
rect 3888 4320 3904 4384
rect 3968 4320 3976 4384
rect 3656 3296 3976 4320
rect 3656 3232 3664 3296
rect 3728 3232 3744 3296
rect 3808 3232 3824 3296
rect 3888 3232 3904 3296
rect 3968 3232 3976 3296
rect 3656 2208 3976 3232
rect 3656 2144 3664 2208
rect 3728 2144 3744 2208
rect 3808 2144 3824 2208
rect 3888 2144 3904 2208
rect 3968 2144 3976 2208
rect 3656 1120 3976 2144
rect 3656 1056 3664 1120
rect 3728 1056 3744 1120
rect 3808 1056 3824 1120
rect 3888 1056 3904 1120
rect 3968 1056 3976 1120
rect 3656 496 3976 1056
rect 4316 19072 4636 19088
rect 4316 19008 4324 19072
rect 4388 19008 4404 19072
rect 4468 19008 4484 19072
rect 4548 19008 4564 19072
rect 4628 19008 4636 19072
rect 4316 17984 4636 19008
rect 4316 17920 4324 17984
rect 4388 17920 4404 17984
rect 4468 17920 4484 17984
rect 4548 17920 4564 17984
rect 4628 17920 4636 17984
rect 4316 16896 4636 17920
rect 4316 16832 4324 16896
rect 4388 16832 4404 16896
rect 4468 16832 4484 16896
rect 4548 16832 4564 16896
rect 4628 16832 4636 16896
rect 4316 15808 4636 16832
rect 4316 15744 4324 15808
rect 4388 15744 4404 15808
rect 4468 15744 4484 15808
rect 4548 15744 4564 15808
rect 4628 15744 4636 15808
rect 4316 14720 4636 15744
rect 4316 14656 4324 14720
rect 4388 14656 4404 14720
rect 4468 14656 4484 14720
rect 4548 14656 4564 14720
rect 4628 14656 4636 14720
rect 4316 13632 4636 14656
rect 4316 13568 4324 13632
rect 4388 13568 4404 13632
rect 4468 13568 4484 13632
rect 4548 13568 4564 13632
rect 4628 13568 4636 13632
rect 4316 12544 4636 13568
rect 4316 12480 4324 12544
rect 4388 12480 4404 12544
rect 4468 12480 4484 12544
rect 4548 12480 4564 12544
rect 4628 12480 4636 12544
rect 4316 11456 4636 12480
rect 4316 11392 4324 11456
rect 4388 11392 4404 11456
rect 4468 11392 4484 11456
rect 4548 11392 4564 11456
rect 4628 11392 4636 11456
rect 4316 10368 4636 11392
rect 4316 10304 4324 10368
rect 4388 10304 4404 10368
rect 4468 10304 4484 10368
rect 4548 10304 4564 10368
rect 4628 10304 4636 10368
rect 4316 9280 4636 10304
rect 4316 9216 4324 9280
rect 4388 9216 4404 9280
rect 4468 9216 4484 9280
rect 4548 9216 4564 9280
rect 4628 9216 4636 9280
rect 4316 8192 4636 9216
rect 4316 8128 4324 8192
rect 4388 8128 4404 8192
rect 4468 8128 4484 8192
rect 4548 8128 4564 8192
rect 4628 8128 4636 8192
rect 4316 7104 4636 8128
rect 4316 7040 4324 7104
rect 4388 7040 4404 7104
rect 4468 7040 4484 7104
rect 4548 7040 4564 7104
rect 4628 7040 4636 7104
rect 4316 6016 4636 7040
rect 4316 5952 4324 6016
rect 4388 5952 4404 6016
rect 4468 5952 4484 6016
rect 4548 5952 4564 6016
rect 4628 5952 4636 6016
rect 4316 4928 4636 5952
rect 4316 4864 4324 4928
rect 4388 4864 4404 4928
rect 4468 4864 4484 4928
rect 4548 4864 4564 4928
rect 4628 4864 4636 4928
rect 4316 3840 4636 4864
rect 4316 3776 4324 3840
rect 4388 3776 4404 3840
rect 4468 3776 4484 3840
rect 4548 3776 4564 3840
rect 4628 3776 4636 3840
rect 4316 2752 4636 3776
rect 4316 2688 4324 2752
rect 4388 2688 4404 2752
rect 4468 2688 4484 2752
rect 4548 2688 4564 2752
rect 4628 2688 4636 2752
rect 4316 1664 4636 2688
rect 4316 1600 4324 1664
rect 4388 1600 4404 1664
rect 4468 1600 4484 1664
rect 4548 1600 4564 1664
rect 4628 1600 4636 1664
rect 4316 576 4636 1600
rect 4316 512 4324 576
rect 4388 512 4404 576
rect 4468 512 4484 576
rect 4548 512 4564 576
rect 4628 512 4636 576
rect 4316 496 4636 512
rect 11430 18528 11750 19088
rect 11430 18464 11438 18528
rect 11502 18464 11518 18528
rect 11582 18464 11598 18528
rect 11662 18464 11678 18528
rect 11742 18464 11750 18528
rect 11430 17440 11750 18464
rect 11430 17376 11438 17440
rect 11502 17376 11518 17440
rect 11582 17376 11598 17440
rect 11662 17376 11678 17440
rect 11742 17376 11750 17440
rect 11430 16352 11750 17376
rect 11430 16288 11438 16352
rect 11502 16288 11518 16352
rect 11582 16288 11598 16352
rect 11662 16288 11678 16352
rect 11742 16288 11750 16352
rect 11430 15264 11750 16288
rect 11430 15200 11438 15264
rect 11502 15200 11518 15264
rect 11582 15200 11598 15264
rect 11662 15200 11678 15264
rect 11742 15200 11750 15264
rect 11430 14176 11750 15200
rect 11430 14112 11438 14176
rect 11502 14112 11518 14176
rect 11582 14112 11598 14176
rect 11662 14112 11678 14176
rect 11742 14112 11750 14176
rect 11430 13088 11750 14112
rect 11430 13024 11438 13088
rect 11502 13024 11518 13088
rect 11582 13024 11598 13088
rect 11662 13024 11678 13088
rect 11742 13024 11750 13088
rect 11430 12000 11750 13024
rect 11430 11936 11438 12000
rect 11502 11936 11518 12000
rect 11582 11936 11598 12000
rect 11662 11936 11678 12000
rect 11742 11936 11750 12000
rect 11430 10912 11750 11936
rect 11430 10848 11438 10912
rect 11502 10848 11518 10912
rect 11582 10848 11598 10912
rect 11662 10848 11678 10912
rect 11742 10848 11750 10912
rect 11430 9824 11750 10848
rect 11430 9760 11438 9824
rect 11502 9760 11518 9824
rect 11582 9760 11598 9824
rect 11662 9760 11678 9824
rect 11742 9760 11750 9824
rect 11430 8736 11750 9760
rect 11430 8672 11438 8736
rect 11502 8672 11518 8736
rect 11582 8672 11598 8736
rect 11662 8672 11678 8736
rect 11742 8672 11750 8736
rect 11430 7648 11750 8672
rect 11430 7584 11438 7648
rect 11502 7584 11518 7648
rect 11582 7584 11598 7648
rect 11662 7584 11678 7648
rect 11742 7584 11750 7648
rect 11430 6560 11750 7584
rect 11430 6496 11438 6560
rect 11502 6496 11518 6560
rect 11582 6496 11598 6560
rect 11662 6496 11678 6560
rect 11742 6496 11750 6560
rect 11430 5472 11750 6496
rect 11430 5408 11438 5472
rect 11502 5408 11518 5472
rect 11582 5408 11598 5472
rect 11662 5408 11678 5472
rect 11742 5408 11750 5472
rect 11430 4384 11750 5408
rect 11430 4320 11438 4384
rect 11502 4320 11518 4384
rect 11582 4320 11598 4384
rect 11662 4320 11678 4384
rect 11742 4320 11750 4384
rect 11430 3296 11750 4320
rect 11430 3232 11438 3296
rect 11502 3232 11518 3296
rect 11582 3232 11598 3296
rect 11662 3232 11678 3296
rect 11742 3232 11750 3296
rect 11430 2208 11750 3232
rect 11430 2144 11438 2208
rect 11502 2144 11518 2208
rect 11582 2144 11598 2208
rect 11662 2144 11678 2208
rect 11742 2144 11750 2208
rect 11430 1120 11750 2144
rect 11430 1056 11438 1120
rect 11502 1056 11518 1120
rect 11582 1056 11598 1120
rect 11662 1056 11678 1120
rect 11742 1056 11750 1120
rect 11430 496 11750 1056
rect 12090 19072 12410 19088
rect 12090 19008 12098 19072
rect 12162 19008 12178 19072
rect 12242 19008 12258 19072
rect 12322 19008 12338 19072
rect 12402 19008 12410 19072
rect 12090 17984 12410 19008
rect 12090 17920 12098 17984
rect 12162 17920 12178 17984
rect 12242 17920 12258 17984
rect 12322 17920 12338 17984
rect 12402 17920 12410 17984
rect 12090 16896 12410 17920
rect 12090 16832 12098 16896
rect 12162 16832 12178 16896
rect 12242 16832 12258 16896
rect 12322 16832 12338 16896
rect 12402 16832 12410 16896
rect 12090 15808 12410 16832
rect 12090 15744 12098 15808
rect 12162 15744 12178 15808
rect 12242 15744 12258 15808
rect 12322 15744 12338 15808
rect 12402 15744 12410 15808
rect 12090 14720 12410 15744
rect 12090 14656 12098 14720
rect 12162 14656 12178 14720
rect 12242 14656 12258 14720
rect 12322 14656 12338 14720
rect 12402 14656 12410 14720
rect 12090 13632 12410 14656
rect 12090 13568 12098 13632
rect 12162 13568 12178 13632
rect 12242 13568 12258 13632
rect 12322 13568 12338 13632
rect 12402 13568 12410 13632
rect 12090 12544 12410 13568
rect 12090 12480 12098 12544
rect 12162 12480 12178 12544
rect 12242 12480 12258 12544
rect 12322 12480 12338 12544
rect 12402 12480 12410 12544
rect 12090 11456 12410 12480
rect 12090 11392 12098 11456
rect 12162 11392 12178 11456
rect 12242 11392 12258 11456
rect 12322 11392 12338 11456
rect 12402 11392 12410 11456
rect 12090 10368 12410 11392
rect 12090 10304 12098 10368
rect 12162 10304 12178 10368
rect 12242 10304 12258 10368
rect 12322 10304 12338 10368
rect 12402 10304 12410 10368
rect 12090 9280 12410 10304
rect 12090 9216 12098 9280
rect 12162 9216 12178 9280
rect 12242 9216 12258 9280
rect 12322 9216 12338 9280
rect 12402 9216 12410 9280
rect 12090 8192 12410 9216
rect 12090 8128 12098 8192
rect 12162 8128 12178 8192
rect 12242 8128 12258 8192
rect 12322 8128 12338 8192
rect 12402 8128 12410 8192
rect 12090 7104 12410 8128
rect 12090 7040 12098 7104
rect 12162 7040 12178 7104
rect 12242 7040 12258 7104
rect 12322 7040 12338 7104
rect 12402 7040 12410 7104
rect 12090 6016 12410 7040
rect 12090 5952 12098 6016
rect 12162 5952 12178 6016
rect 12242 5952 12258 6016
rect 12322 5952 12338 6016
rect 12402 5952 12410 6016
rect 12090 4928 12410 5952
rect 12090 4864 12098 4928
rect 12162 4864 12178 4928
rect 12242 4864 12258 4928
rect 12322 4864 12338 4928
rect 12402 4864 12410 4928
rect 12090 3840 12410 4864
rect 12090 3776 12098 3840
rect 12162 3776 12178 3840
rect 12242 3776 12258 3840
rect 12322 3776 12338 3840
rect 12402 3776 12410 3840
rect 12090 2752 12410 3776
rect 12090 2688 12098 2752
rect 12162 2688 12178 2752
rect 12242 2688 12258 2752
rect 12322 2688 12338 2752
rect 12402 2688 12410 2752
rect 12090 1664 12410 2688
rect 12090 1600 12098 1664
rect 12162 1600 12178 1664
rect 12242 1600 12258 1664
rect 12322 1600 12338 1664
rect 12402 1600 12410 1664
rect 12090 576 12410 1600
rect 12090 512 12098 576
rect 12162 512 12178 576
rect 12242 512 12258 576
rect 12322 512 12338 576
rect 12402 512 12410 576
rect 12090 496 12410 512
rect 19204 18528 19524 19088
rect 19204 18464 19212 18528
rect 19276 18464 19292 18528
rect 19356 18464 19372 18528
rect 19436 18464 19452 18528
rect 19516 18464 19524 18528
rect 19204 17440 19524 18464
rect 19204 17376 19212 17440
rect 19276 17376 19292 17440
rect 19356 17376 19372 17440
rect 19436 17376 19452 17440
rect 19516 17376 19524 17440
rect 19204 16352 19524 17376
rect 19204 16288 19212 16352
rect 19276 16288 19292 16352
rect 19356 16288 19372 16352
rect 19436 16288 19452 16352
rect 19516 16288 19524 16352
rect 19204 15264 19524 16288
rect 19204 15200 19212 15264
rect 19276 15200 19292 15264
rect 19356 15200 19372 15264
rect 19436 15200 19452 15264
rect 19516 15200 19524 15264
rect 19204 14176 19524 15200
rect 19204 14112 19212 14176
rect 19276 14112 19292 14176
rect 19356 14112 19372 14176
rect 19436 14112 19452 14176
rect 19516 14112 19524 14176
rect 19204 13088 19524 14112
rect 19204 13024 19212 13088
rect 19276 13024 19292 13088
rect 19356 13024 19372 13088
rect 19436 13024 19452 13088
rect 19516 13024 19524 13088
rect 19204 12000 19524 13024
rect 19204 11936 19212 12000
rect 19276 11936 19292 12000
rect 19356 11936 19372 12000
rect 19436 11936 19452 12000
rect 19516 11936 19524 12000
rect 19204 10912 19524 11936
rect 19204 10848 19212 10912
rect 19276 10848 19292 10912
rect 19356 10848 19372 10912
rect 19436 10848 19452 10912
rect 19516 10848 19524 10912
rect 19204 9824 19524 10848
rect 19204 9760 19212 9824
rect 19276 9760 19292 9824
rect 19356 9760 19372 9824
rect 19436 9760 19452 9824
rect 19516 9760 19524 9824
rect 19204 8736 19524 9760
rect 19204 8672 19212 8736
rect 19276 8672 19292 8736
rect 19356 8672 19372 8736
rect 19436 8672 19452 8736
rect 19516 8672 19524 8736
rect 19204 7648 19524 8672
rect 19204 7584 19212 7648
rect 19276 7584 19292 7648
rect 19356 7584 19372 7648
rect 19436 7584 19452 7648
rect 19516 7584 19524 7648
rect 19204 6560 19524 7584
rect 19204 6496 19212 6560
rect 19276 6496 19292 6560
rect 19356 6496 19372 6560
rect 19436 6496 19452 6560
rect 19516 6496 19524 6560
rect 19204 5472 19524 6496
rect 19204 5408 19212 5472
rect 19276 5408 19292 5472
rect 19356 5408 19372 5472
rect 19436 5408 19452 5472
rect 19516 5408 19524 5472
rect 19204 4384 19524 5408
rect 19204 4320 19212 4384
rect 19276 4320 19292 4384
rect 19356 4320 19372 4384
rect 19436 4320 19452 4384
rect 19516 4320 19524 4384
rect 19204 3296 19524 4320
rect 19204 3232 19212 3296
rect 19276 3232 19292 3296
rect 19356 3232 19372 3296
rect 19436 3232 19452 3296
rect 19516 3232 19524 3296
rect 19204 2208 19524 3232
rect 19204 2144 19212 2208
rect 19276 2144 19292 2208
rect 19356 2144 19372 2208
rect 19436 2144 19452 2208
rect 19516 2144 19524 2208
rect 19204 1120 19524 2144
rect 19204 1056 19212 1120
rect 19276 1056 19292 1120
rect 19356 1056 19372 1120
rect 19436 1056 19452 1120
rect 19516 1056 19524 1120
rect 19204 496 19524 1056
rect 19864 19072 20184 19088
rect 19864 19008 19872 19072
rect 19936 19008 19952 19072
rect 20016 19008 20032 19072
rect 20096 19008 20112 19072
rect 20176 19008 20184 19072
rect 19864 17984 20184 19008
rect 19864 17920 19872 17984
rect 19936 17920 19952 17984
rect 20016 17920 20032 17984
rect 20096 17920 20112 17984
rect 20176 17920 20184 17984
rect 19864 16896 20184 17920
rect 19864 16832 19872 16896
rect 19936 16832 19952 16896
rect 20016 16832 20032 16896
rect 20096 16832 20112 16896
rect 20176 16832 20184 16896
rect 19864 15808 20184 16832
rect 19864 15744 19872 15808
rect 19936 15744 19952 15808
rect 20016 15744 20032 15808
rect 20096 15744 20112 15808
rect 20176 15744 20184 15808
rect 19864 14720 20184 15744
rect 19864 14656 19872 14720
rect 19936 14656 19952 14720
rect 20016 14656 20032 14720
rect 20096 14656 20112 14720
rect 20176 14656 20184 14720
rect 19864 13632 20184 14656
rect 19864 13568 19872 13632
rect 19936 13568 19952 13632
rect 20016 13568 20032 13632
rect 20096 13568 20112 13632
rect 20176 13568 20184 13632
rect 19864 12544 20184 13568
rect 19864 12480 19872 12544
rect 19936 12480 19952 12544
rect 20016 12480 20032 12544
rect 20096 12480 20112 12544
rect 20176 12480 20184 12544
rect 19864 11456 20184 12480
rect 19864 11392 19872 11456
rect 19936 11392 19952 11456
rect 20016 11392 20032 11456
rect 20096 11392 20112 11456
rect 20176 11392 20184 11456
rect 19864 10368 20184 11392
rect 19864 10304 19872 10368
rect 19936 10304 19952 10368
rect 20016 10304 20032 10368
rect 20096 10304 20112 10368
rect 20176 10304 20184 10368
rect 19864 9280 20184 10304
rect 19864 9216 19872 9280
rect 19936 9216 19952 9280
rect 20016 9216 20032 9280
rect 20096 9216 20112 9280
rect 20176 9216 20184 9280
rect 19864 8192 20184 9216
rect 19864 8128 19872 8192
rect 19936 8128 19952 8192
rect 20016 8128 20032 8192
rect 20096 8128 20112 8192
rect 20176 8128 20184 8192
rect 19864 7104 20184 8128
rect 19864 7040 19872 7104
rect 19936 7040 19952 7104
rect 20016 7040 20032 7104
rect 20096 7040 20112 7104
rect 20176 7040 20184 7104
rect 19864 6016 20184 7040
rect 19864 5952 19872 6016
rect 19936 5952 19952 6016
rect 20016 5952 20032 6016
rect 20096 5952 20112 6016
rect 20176 5952 20184 6016
rect 19864 4928 20184 5952
rect 19864 4864 19872 4928
rect 19936 4864 19952 4928
rect 20016 4864 20032 4928
rect 20096 4864 20112 4928
rect 20176 4864 20184 4928
rect 19864 3840 20184 4864
rect 19864 3776 19872 3840
rect 19936 3776 19952 3840
rect 20016 3776 20032 3840
rect 20096 3776 20112 3840
rect 20176 3776 20184 3840
rect 19864 2752 20184 3776
rect 19864 2688 19872 2752
rect 19936 2688 19952 2752
rect 20016 2688 20032 2752
rect 20096 2688 20112 2752
rect 20176 2688 20184 2752
rect 19864 1664 20184 2688
rect 19864 1600 19872 1664
rect 19936 1600 19952 1664
rect 20016 1600 20032 1664
rect 20096 1600 20112 1664
rect 20176 1600 20184 1664
rect 19864 576 20184 1600
rect 19864 512 19872 576
rect 19936 512 19952 576
rect 20016 512 20032 576
rect 20096 512 20112 576
rect 20176 512 20184 576
rect 19864 496 20184 512
rect 26978 18528 27298 19088
rect 26978 18464 26986 18528
rect 27050 18464 27066 18528
rect 27130 18464 27146 18528
rect 27210 18464 27226 18528
rect 27290 18464 27298 18528
rect 26978 17440 27298 18464
rect 26978 17376 26986 17440
rect 27050 17376 27066 17440
rect 27130 17376 27146 17440
rect 27210 17376 27226 17440
rect 27290 17376 27298 17440
rect 26978 16352 27298 17376
rect 26978 16288 26986 16352
rect 27050 16288 27066 16352
rect 27130 16288 27146 16352
rect 27210 16288 27226 16352
rect 27290 16288 27298 16352
rect 26978 15264 27298 16288
rect 26978 15200 26986 15264
rect 27050 15200 27066 15264
rect 27130 15200 27146 15264
rect 27210 15200 27226 15264
rect 27290 15200 27298 15264
rect 26978 14176 27298 15200
rect 26978 14112 26986 14176
rect 27050 14112 27066 14176
rect 27130 14112 27146 14176
rect 27210 14112 27226 14176
rect 27290 14112 27298 14176
rect 26978 13088 27298 14112
rect 26978 13024 26986 13088
rect 27050 13024 27066 13088
rect 27130 13024 27146 13088
rect 27210 13024 27226 13088
rect 27290 13024 27298 13088
rect 26978 12000 27298 13024
rect 26978 11936 26986 12000
rect 27050 11936 27066 12000
rect 27130 11936 27146 12000
rect 27210 11936 27226 12000
rect 27290 11936 27298 12000
rect 26978 10912 27298 11936
rect 26978 10848 26986 10912
rect 27050 10848 27066 10912
rect 27130 10848 27146 10912
rect 27210 10848 27226 10912
rect 27290 10848 27298 10912
rect 26978 9824 27298 10848
rect 26978 9760 26986 9824
rect 27050 9760 27066 9824
rect 27130 9760 27146 9824
rect 27210 9760 27226 9824
rect 27290 9760 27298 9824
rect 26978 8736 27298 9760
rect 26978 8672 26986 8736
rect 27050 8672 27066 8736
rect 27130 8672 27146 8736
rect 27210 8672 27226 8736
rect 27290 8672 27298 8736
rect 26978 7648 27298 8672
rect 26978 7584 26986 7648
rect 27050 7584 27066 7648
rect 27130 7584 27146 7648
rect 27210 7584 27226 7648
rect 27290 7584 27298 7648
rect 26978 6560 27298 7584
rect 26978 6496 26986 6560
rect 27050 6496 27066 6560
rect 27130 6496 27146 6560
rect 27210 6496 27226 6560
rect 27290 6496 27298 6560
rect 26978 5472 27298 6496
rect 26978 5408 26986 5472
rect 27050 5408 27066 5472
rect 27130 5408 27146 5472
rect 27210 5408 27226 5472
rect 27290 5408 27298 5472
rect 26978 4384 27298 5408
rect 26978 4320 26986 4384
rect 27050 4320 27066 4384
rect 27130 4320 27146 4384
rect 27210 4320 27226 4384
rect 27290 4320 27298 4384
rect 26978 3296 27298 4320
rect 26978 3232 26986 3296
rect 27050 3232 27066 3296
rect 27130 3232 27146 3296
rect 27210 3232 27226 3296
rect 27290 3232 27298 3296
rect 26978 2208 27298 3232
rect 26978 2144 26986 2208
rect 27050 2144 27066 2208
rect 27130 2144 27146 2208
rect 27210 2144 27226 2208
rect 27290 2144 27298 2208
rect 26978 1120 27298 2144
rect 26978 1056 26986 1120
rect 27050 1056 27066 1120
rect 27130 1056 27146 1120
rect 27210 1056 27226 1120
rect 27290 1056 27298 1120
rect 26978 496 27298 1056
rect 27638 19072 27958 19088
rect 27638 19008 27646 19072
rect 27710 19008 27726 19072
rect 27790 19008 27806 19072
rect 27870 19008 27886 19072
rect 27950 19008 27958 19072
rect 27638 17984 27958 19008
rect 27638 17920 27646 17984
rect 27710 17920 27726 17984
rect 27790 17920 27806 17984
rect 27870 17920 27886 17984
rect 27950 17920 27958 17984
rect 27638 16896 27958 17920
rect 27638 16832 27646 16896
rect 27710 16832 27726 16896
rect 27790 16832 27806 16896
rect 27870 16832 27886 16896
rect 27950 16832 27958 16896
rect 27638 15808 27958 16832
rect 27638 15744 27646 15808
rect 27710 15744 27726 15808
rect 27790 15744 27806 15808
rect 27870 15744 27886 15808
rect 27950 15744 27958 15808
rect 27638 14720 27958 15744
rect 27638 14656 27646 14720
rect 27710 14656 27726 14720
rect 27790 14656 27806 14720
rect 27870 14656 27886 14720
rect 27950 14656 27958 14720
rect 27638 13632 27958 14656
rect 27638 13568 27646 13632
rect 27710 13568 27726 13632
rect 27790 13568 27806 13632
rect 27870 13568 27886 13632
rect 27950 13568 27958 13632
rect 27638 12544 27958 13568
rect 27638 12480 27646 12544
rect 27710 12480 27726 12544
rect 27790 12480 27806 12544
rect 27870 12480 27886 12544
rect 27950 12480 27958 12544
rect 27638 11456 27958 12480
rect 27638 11392 27646 11456
rect 27710 11392 27726 11456
rect 27790 11392 27806 11456
rect 27870 11392 27886 11456
rect 27950 11392 27958 11456
rect 27638 10368 27958 11392
rect 27638 10304 27646 10368
rect 27710 10304 27726 10368
rect 27790 10304 27806 10368
rect 27870 10304 27886 10368
rect 27950 10304 27958 10368
rect 27638 9280 27958 10304
rect 27638 9216 27646 9280
rect 27710 9216 27726 9280
rect 27790 9216 27806 9280
rect 27870 9216 27886 9280
rect 27950 9216 27958 9280
rect 27638 8192 27958 9216
rect 27638 8128 27646 8192
rect 27710 8128 27726 8192
rect 27790 8128 27806 8192
rect 27870 8128 27886 8192
rect 27950 8128 27958 8192
rect 27638 7104 27958 8128
rect 27638 7040 27646 7104
rect 27710 7040 27726 7104
rect 27790 7040 27806 7104
rect 27870 7040 27886 7104
rect 27950 7040 27958 7104
rect 27638 6016 27958 7040
rect 27638 5952 27646 6016
rect 27710 5952 27726 6016
rect 27790 5952 27806 6016
rect 27870 5952 27886 6016
rect 27950 5952 27958 6016
rect 27638 4928 27958 5952
rect 27638 4864 27646 4928
rect 27710 4864 27726 4928
rect 27790 4864 27806 4928
rect 27870 4864 27886 4928
rect 27950 4864 27958 4928
rect 27638 3840 27958 4864
rect 27638 3776 27646 3840
rect 27710 3776 27726 3840
rect 27790 3776 27806 3840
rect 27870 3776 27886 3840
rect 27950 3776 27958 3840
rect 27638 2752 27958 3776
rect 27638 2688 27646 2752
rect 27710 2688 27726 2752
rect 27790 2688 27806 2752
rect 27870 2688 27886 2752
rect 27950 2688 27958 2752
rect 27638 1664 27958 2688
rect 27638 1600 27646 1664
rect 27710 1600 27726 1664
rect 27790 1600 27806 1664
rect 27870 1600 27886 1664
rect 27950 1600 27958 1664
rect 27638 576 27958 1600
rect 27638 512 27646 576
rect 27710 512 27726 576
rect 27790 512 27806 576
rect 27870 512 27886 576
rect 27950 512 27958 576
rect 27638 496 27958 512
use sky130_fd_sc_hd__inv_2  _033_
timestamp 18001
transform -1 0 14996 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _034_
timestamp 18001
transform -1 0 15640 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _035_
timestamp 18001
transform 1 0 18124 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _036_
timestamp 18001
transform 1 0 14720 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _037_
timestamp 18001
transform -1 0 17296 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__or4_2  _038_
timestamp 18001
transform -1 0 16836 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__o22ai_1  _039_
timestamp 18001
transform 1 0 14076 0 -1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _040_
timestamp 18001
transform 1 0 14628 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__o41a_2  _041_
timestamp 18001
transform 1 0 16100 0 -1 16864
box -38 -48 958 592
use sky130_fd_sc_hd__o21a_1  _042_
timestamp 18001
transform -1 0 17480 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _043_
timestamp 18001
transform 1 0 17388 0 1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _044_
timestamp 18001
transform -1 0 18216 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _045_
timestamp 18001
transform -1 0 17112 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _046_
timestamp 18001
transform -1 0 17664 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _047_
timestamp 18001
transform -1 0 17204 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _048_
timestamp 18001
transform -1 0 17388 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _049_
timestamp 18001
transform -1 0 18584 0 1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _050_
timestamp 18001
transform 1 0 17112 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__and3_2  _051_
timestamp 18001
transform -1 0 16836 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _052_
timestamp 18001
transform -1 0 16008 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _053_
timestamp 18001
transform -1 0 17572 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _054_
timestamp 18001
transform -1 0 14260 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__o2111a_1  _055_
timestamp 18001
transform 1 0 14536 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _056_
timestamp 18001
transform 1 0 13524 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _057_
timestamp 18001
transform -1 0 14720 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _058_
timestamp 18001
transform -1 0 13340 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _059_
timestamp 18001
transform -1 0 16008 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_1  _060_
timestamp 18001
transform 1 0 12328 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _061_
timestamp 18001
transform -1 0 13432 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__nand4_1  _062_
timestamp 18001
transform 1 0 13524 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _063_
timestamp 18001
transform 1 0 14904 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _064_
timestamp 18001
transform 1 0 14536 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _065_
timestamp 18001
transform 1 0 16100 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__dfrtp_1  _066_
timestamp 18001
transform -1 0 19320 0 -1 17952
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _067_
timestamp 18001
transform 1 0 16468 0 -1 14688
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _068_
timestamp 18001
transform 1 0 17572 0 -1 15776
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _069_
timestamp 18001
transform -1 0 19228 0 -1 16864
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _070_
timestamp 18001
transform 1 0 12236 0 -1 17952
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _071_
timestamp 18001
transform 1 0 12236 0 -1 15776
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _072_
timestamp 18001
transform 1 0 12696 0 -1 14688
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _073_
timestamp 18001
transform -1 0 15364 0 1 13600
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _074_
timestamp 18001
transform 1 0 13524 0 1 17952
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _075_
timestamp 18001
transform 1 0 14996 0 1 16864
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _076_
timestamp 18001
transform 1 0 15456 0 1 17952
box -38 -48 1970 592
use sky130_fd_sc_hd__buf_2  _098_
timestamp 18001
transform 1 0 17756 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _099_
timestamp 18001
transform 1 0 17848 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _100_
timestamp 18001
transform -1 0 14996 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp 18001
transform -1 0 16836 0 1 15776
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_clk
timestamp 18001
transform -1 0 14536 0 -1 16864
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_clk
timestamp 18001
transform 1 0 19228 0 -1 16864
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_4  clkload0
timestamp 18001
transform 1 0 12696 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout3
timestamp 18001
transform 1 0 18216 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout4
timestamp 18001
transform 1 0 18308 0 -1 14688
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3
timestamp 1636986456
transform 1 0 828 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 1636986456
transform 1 0 1932 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27
timestamp 18001
transform 1 0 3036 0 1 544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1636986456
transform 1 0 3220 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1636986456
transform 1 0 4324 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53
timestamp 18001
transform 1 0 5428 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1636986456
transform 1 0 5796 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_69
timestamp 18001
transform 1 0 6900 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_75
timestamp 18001
transform 1 0 7452 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83
timestamp 18001
transform 1 0 8188 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_85
timestamp 18001
transform 1 0 8372 0 1 544
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96
timestamp 1636986456
transform 1 0 9384 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_108
timestamp 18001
transform 1 0 10488 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_113
timestamp 18001
transform 1 0 10948 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_124
timestamp 18001
transform 1 0 11960 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_131
timestamp 18001
transform 1 0 12604 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_138
timestamp 18001
transform 1 0 13248 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_141
timestamp 18001
transform 1 0 13524 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_145
timestamp 18001
transform 1 0 13892 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_152
timestamp 18001
transform 1 0 14536 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_159
timestamp 18001
transform 1 0 15180 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_166
timestamp 18001
transform 1 0 15824 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_169
timestamp 18001
transform 1 0 16100 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_180
timestamp 18001
transform 1 0 17112 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_187
timestamp 18001
transform 1 0 17756 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_194
timestamp 18001
transform 1 0 18400 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_197
timestamp 18001
transform 1 0 18676 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_201
timestamp 18001
transform 1 0 19044 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_209
timestamp 18001
transform 1 0 19780 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_215
timestamp 18001
transform 1 0 20332 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_223
timestamp 18001
transform 1 0 21068 0 1 544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_225
timestamp 1636986456
transform 1 0 21252 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_237
timestamp 1636986456
transform 1 0 22356 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp 18001
transform 1 0 23460 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_253
timestamp 1636986456
transform 1 0 23828 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_265
timestamp 1636986456
transform 1 0 24932 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_277
timestamp 18001
transform 1 0 26036 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_281
timestamp 1636986456
transform 1 0 26404 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_293
timestamp 1636986456
transform 1 0 27508 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_305
timestamp 18001
transform 1 0 28612 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_309
timestamp 1636986456
transform 1 0 28980 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_321
timestamp 18001
transform 1 0 30084 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_329
timestamp 18001
transform 1 0 30820 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1636986456
transform 1 0 828 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1636986456
transform 1 0 1932 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1636986456
transform 1 0 3036 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1636986456
transform 1 0 4140 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 18001
transform 1 0 5244 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 18001
transform 1 0 5612 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1636986456
transform 1 0 5796 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1636986456
transform 1 0 6900 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1636986456
transform 1 0 8004 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1636986456
transform 1 0 9108 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 18001
transform 1 0 10212 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 18001
transform 1 0 10764 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1636986456
transform 1 0 10948 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1636986456
transform 1 0 12052 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1636986456
transform 1 0 13156 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1636986456
transform 1 0 14260 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 18001
transform 1 0 15364 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 18001
transform 1 0 15916 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1636986456
transform 1 0 16100 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_181
timestamp 1636986456
transform 1 0 17204 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_193
timestamp 1636986456
transform 1 0 18308 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_205
timestamp 1636986456
transform 1 0 19412 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp 18001
transform 1 0 20516 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 18001
transform 1 0 21068 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1636986456
transform 1 0 21252 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_237
timestamp 1636986456
transform 1 0 22356 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_249
timestamp 1636986456
transform 1 0 23460 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_261
timestamp 1636986456
transform 1 0 24564 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp 18001
transform 1 0 25668 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 18001
transform 1 0 26220 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_281
timestamp 1636986456
transform 1 0 26404 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_293
timestamp 1636986456
transform 1 0 27508 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_305
timestamp 1636986456
transform 1 0 28612 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_317
timestamp 1636986456
transform 1 0 29716 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_329
timestamp 18001
transform 1 0 30820 0 -1 1632
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1636986456
transform 1 0 828 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1636986456
transform 1 0 1932 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 18001
transform 1 0 3036 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1636986456
transform 1 0 3220 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1636986456
transform 1 0 4324 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1636986456
transform 1 0 5428 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1636986456
transform 1 0 6532 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 18001
transform 1 0 7636 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 18001
transform 1 0 8188 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1636986456
transform 1 0 8372 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1636986456
transform 1 0 9476 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1636986456
transform 1 0 10580 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1636986456
transform 1 0 11684 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 18001
transform 1 0 12788 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 18001
transform 1 0 13340 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1636986456
transform 1 0 13524 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1636986456
transform 1 0 14628 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1636986456
transform 1 0 15732 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1636986456
transform 1 0 16836 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 18001
transform 1 0 17940 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 18001
transform 1 0 18492 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1636986456
transform 1 0 18676 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1636986456
transform 1 0 19780 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_221
timestamp 1636986456
transform 1 0 20884 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_233
timestamp 1636986456
transform 1 0 21988 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 18001
transform 1 0 23092 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 18001
transform 1 0 23644 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1636986456
transform 1 0 23828 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_265
timestamp 1636986456
transform 1 0 24932 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_277
timestamp 1636986456
transform 1 0 26036 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_289
timestamp 1636986456
transform 1 0 27140 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp 18001
transform 1 0 28244 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 18001
transform 1 0 28796 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1636986456
transform 1 0 28980 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_321
timestamp 18001
transform 1 0 30084 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_329
timestamp 18001
transform 1 0 30820 0 1 1632
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1636986456
transform 1 0 828 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1636986456
transform 1 0 1932 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1636986456
transform 1 0 3036 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1636986456
transform 1 0 4140 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 18001
transform 1 0 5244 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 18001
transform 1 0 5612 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1636986456
transform 1 0 5796 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1636986456
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1636986456
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1636986456
transform 1 0 9108 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 18001
transform 1 0 10212 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 18001
transform 1 0 10764 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1636986456
transform 1 0 10948 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1636986456
transform 1 0 12052 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1636986456
transform 1 0 13156 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1636986456
transform 1 0 14260 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 18001
transform 1 0 15364 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 18001
transform 1 0 15916 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1636986456
transform 1 0 16100 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1636986456
transform 1 0 17204 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1636986456
transform 1 0 18308 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1636986456
transform 1 0 19412 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 18001
transform 1 0 20516 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 18001
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1636986456
transform 1 0 21252 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1636986456
transform 1 0 22356 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_249
timestamp 1636986456
transform 1 0 23460 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_261
timestamp 1636986456
transform 1 0 24564 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 18001
transform 1 0 25668 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 18001
transform 1 0 26220 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1636986456
transform 1 0 26404 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1636986456
transform 1 0 27508 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_305
timestamp 1636986456
transform 1 0 28612 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_317
timestamp 1636986456
transform 1 0 29716 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_329
timestamp 18001
transform 1 0 30820 0 -1 2720
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1636986456
transform 1 0 828 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1636986456
transform 1 0 1932 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 18001
transform 1 0 3036 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1636986456
transform 1 0 3220 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1636986456
transform 1 0 4324 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1636986456
transform 1 0 5428 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1636986456
transform 1 0 6532 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 18001
transform 1 0 7636 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 18001
transform 1 0 8188 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1636986456
transform 1 0 8372 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1636986456
transform 1 0 9476 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1636986456
transform 1 0 10580 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1636986456
transform 1 0 11684 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 18001
transform 1 0 12788 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 18001
transform 1 0 13340 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1636986456
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1636986456
transform 1 0 14628 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1636986456
transform 1 0 15732 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1636986456
transform 1 0 16836 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 18001
transform 1 0 17940 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 18001
transform 1 0 18492 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1636986456
transform 1 0 18676 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1636986456
transform 1 0 19780 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_221
timestamp 1636986456
transform 1 0 20884 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_233
timestamp 1636986456
transform 1 0 21988 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 18001
transform 1 0 23092 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 18001
transform 1 0 23644 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1636986456
transform 1 0 23828 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1636986456
transform 1 0 24932 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_277
timestamp 1636986456
transform 1 0 26036 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_289
timestamp 1636986456
transform 1 0 27140 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 18001
transform 1 0 28244 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 18001
transform 1 0 28796 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1636986456
transform 1 0 28980 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_321
timestamp 18001
transform 1 0 30084 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_329
timestamp 18001
transform 1 0 30820 0 1 2720
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1636986456
transform 1 0 828 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1636986456
transform 1 0 1932 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1636986456
transform 1 0 3036 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1636986456
transform 1 0 4140 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 18001
transform 1 0 5244 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 18001
transform 1 0 5612 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1636986456
transform 1 0 5796 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1636986456
transform 1 0 6900 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1636986456
transform 1 0 8004 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1636986456
transform 1 0 9108 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 18001
transform 1 0 10212 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 18001
transform 1 0 10764 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1636986456
transform 1 0 10948 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1636986456
transform 1 0 12052 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1636986456
transform 1 0 13156 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1636986456
transform 1 0 14260 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 18001
transform 1 0 15364 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 18001
transform 1 0 15916 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1636986456
transform 1 0 16100 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1636986456
transform 1 0 17204 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1636986456
transform 1 0 18308 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1636986456
transform 1 0 19412 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 18001
transform 1 0 20516 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 18001
transform 1 0 21068 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1636986456
transform 1 0 21252 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1636986456
transform 1 0 22356 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_249
timestamp 1636986456
transform 1 0 23460 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_261
timestamp 1636986456
transform 1 0 24564 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 18001
transform 1 0 25668 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 18001
transform 1 0 26220 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1636986456
transform 1 0 26404 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_293
timestamp 1636986456
transform 1 0 27508 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_305
timestamp 1636986456
transform 1 0 28612 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_317
timestamp 1636986456
transform 1 0 29716 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_329
timestamp 18001
transform 1 0 30820 0 -1 3808
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1636986456
transform 1 0 828 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1636986456
transform 1 0 1932 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 18001
transform 1 0 3036 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1636986456
transform 1 0 3220 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1636986456
transform 1 0 4324 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1636986456
transform 1 0 5428 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1636986456
transform 1 0 6532 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 18001
transform 1 0 7636 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 18001
transform 1 0 8188 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1636986456
transform 1 0 8372 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1636986456
transform 1 0 9476 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1636986456
transform 1 0 10580 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1636986456
transform 1 0 11684 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 18001
transform 1 0 12788 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 18001
transform 1 0 13340 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1636986456
transform 1 0 13524 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1636986456
transform 1 0 14628 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1636986456
transform 1 0 15732 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1636986456
transform 1 0 16836 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 18001
transform 1 0 17940 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 18001
transform 1 0 18492 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1636986456
transform 1 0 18676 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1636986456
transform 1 0 19780 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_221
timestamp 1636986456
transform 1 0 20884 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_233
timestamp 1636986456
transform 1 0 21988 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 18001
transform 1 0 23092 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 18001
transform 1 0 23644 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1636986456
transform 1 0 23828 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1636986456
transform 1 0 24932 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_277
timestamp 1636986456
transform 1 0 26036 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_289
timestamp 1636986456
transform 1 0 27140 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 18001
transform 1 0 28244 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 18001
transform 1 0 28796 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1636986456
transform 1 0 28980 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_321
timestamp 18001
transform 1 0 30084 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_329
timestamp 18001
transform 1 0 30820 0 1 3808
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1636986456
transform 1 0 828 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1636986456
transform 1 0 1932 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1636986456
transform 1 0 3036 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1636986456
transform 1 0 4140 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 18001
transform 1 0 5244 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 18001
transform 1 0 5612 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1636986456
transform 1 0 5796 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1636986456
transform 1 0 6900 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1636986456
transform 1 0 8004 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1636986456
transform 1 0 9108 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 18001
transform 1 0 10212 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 18001
transform 1 0 10764 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1636986456
transform 1 0 10948 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1636986456
transform 1 0 12052 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1636986456
transform 1 0 13156 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1636986456
transform 1 0 14260 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 18001
transform 1 0 15364 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 18001
transform 1 0 15916 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1636986456
transform 1 0 16100 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1636986456
transform 1 0 17204 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1636986456
transform 1 0 18308 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1636986456
transform 1 0 19412 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 18001
transform 1 0 20516 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 18001
transform 1 0 21068 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1636986456
transform 1 0 21252 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1636986456
transform 1 0 22356 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_249
timestamp 1636986456
transform 1 0 23460 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_261
timestamp 1636986456
transform 1 0 24564 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 18001
transform 1 0 25668 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 18001
transform 1 0 26220 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1636986456
transform 1 0 26404 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_293
timestamp 1636986456
transform 1 0 27508 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_305
timestamp 1636986456
transform 1 0 28612 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_317
timestamp 1636986456
transform 1 0 29716 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_329
timestamp 18001
transform 1 0 30820 0 -1 4896
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1636986456
transform 1 0 828 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1636986456
transform 1 0 1932 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 18001
transform 1 0 3036 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1636986456
transform 1 0 3220 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1636986456
transform 1 0 4324 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1636986456
transform 1 0 5428 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1636986456
transform 1 0 6532 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 18001
transform 1 0 7636 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 18001
transform 1 0 8188 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1636986456
transform 1 0 8372 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1636986456
transform 1 0 9476 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1636986456
transform 1 0 10580 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1636986456
transform 1 0 11684 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 18001
transform 1 0 12788 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 18001
transform 1 0 13340 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1636986456
transform 1 0 13524 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1636986456
transform 1 0 14628 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1636986456
transform 1 0 15732 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1636986456
transform 1 0 16836 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 18001
transform 1 0 17940 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 18001
transform 1 0 18492 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1636986456
transform 1 0 18676 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1636986456
transform 1 0 19780 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_221
timestamp 1636986456
transform 1 0 20884 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_233
timestamp 1636986456
transform 1 0 21988 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 18001
transform 1 0 23092 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 18001
transform 1 0 23644 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1636986456
transform 1 0 23828 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1636986456
transform 1 0 24932 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_277
timestamp 1636986456
transform 1 0 26036 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_289
timestamp 1636986456
transform 1 0 27140 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 18001
transform 1 0 28244 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 18001
transform 1 0 28796 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1636986456
transform 1 0 28980 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_321
timestamp 18001
transform 1 0 30084 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_329
timestamp 18001
transform 1 0 30820 0 1 4896
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1636986456
transform 1 0 828 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1636986456
transform 1 0 1932 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1636986456
transform 1 0 3036 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1636986456
transform 1 0 4140 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 18001
transform 1 0 5244 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 18001
transform 1 0 5612 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1636986456
transform 1 0 5796 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1636986456
transform 1 0 6900 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1636986456
transform 1 0 8004 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1636986456
transform 1 0 9108 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 18001
transform 1 0 10212 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 18001
transform 1 0 10764 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1636986456
transform 1 0 10948 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1636986456
transform 1 0 12052 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1636986456
transform 1 0 13156 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1636986456
transform 1 0 14260 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 18001
transform 1 0 15364 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 18001
transform 1 0 15916 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1636986456
transform 1 0 16100 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1636986456
transform 1 0 17204 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_193
timestamp 1636986456
transform 1 0 18308 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_205
timestamp 1636986456
transform 1 0 19412 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 18001
transform 1 0 20516 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 18001
transform 1 0 21068 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_225
timestamp 1636986456
transform 1 0 21252 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_237
timestamp 1636986456
transform 1 0 22356 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_249
timestamp 1636986456
transform 1 0 23460 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_261
timestamp 1636986456
transform 1 0 24564 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 18001
transform 1 0 25668 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 18001
transform 1 0 26220 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1636986456
transform 1 0 26404 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1636986456
transform 1 0 27508 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_305
timestamp 1636986456
transform 1 0 28612 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_317
timestamp 1636986456
transform 1 0 29716 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_329
timestamp 18001
transform 1 0 30820 0 -1 5984
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1636986456
transform 1 0 828 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1636986456
transform 1 0 1932 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 18001
transform 1 0 3036 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1636986456
transform 1 0 3220 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1636986456
transform 1 0 4324 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1636986456
transform 1 0 5428 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1636986456
transform 1 0 6532 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 18001
transform 1 0 7636 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 18001
transform 1 0 8188 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1636986456
transform 1 0 8372 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1636986456
transform 1 0 9476 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1636986456
transform 1 0 10580 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1636986456
transform 1 0 11684 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 18001
transform 1 0 12788 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 18001
transform 1 0 13340 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1636986456
transform 1 0 13524 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1636986456
transform 1 0 14628 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1636986456
transform 1 0 15732 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1636986456
transform 1 0 16836 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 18001
transform 1 0 17940 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 18001
transform 1 0 18492 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1636986456
transform 1 0 18676 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_209
timestamp 1636986456
transform 1 0 19780 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_221
timestamp 1636986456
transform 1 0 20884 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_233
timestamp 1636986456
transform 1 0 21988 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 18001
transform 1 0 23092 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 18001
transform 1 0 23644 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1636986456
transform 1 0 23828 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_265
timestamp 1636986456
transform 1 0 24932 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_277
timestamp 1636986456
transform 1 0 26036 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_289
timestamp 1636986456
transform 1 0 27140 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 18001
transform 1 0 28244 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 18001
transform 1 0 28796 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_309
timestamp 1636986456
transform 1 0 28980 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_321
timestamp 18001
transform 1 0 30084 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_329
timestamp 18001
transform 1 0 30820 0 1 5984
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1636986456
transform 1 0 828 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1636986456
transform 1 0 1932 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1636986456
transform 1 0 3036 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1636986456
transform 1 0 4140 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 18001
transform 1 0 5244 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 18001
transform 1 0 5612 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1636986456
transform 1 0 5796 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1636986456
transform 1 0 6900 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1636986456
transform 1 0 8004 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1636986456
transform 1 0 9108 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 18001
transform 1 0 10212 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 18001
transform 1 0 10764 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1636986456
transform 1 0 10948 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1636986456
transform 1 0 12052 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1636986456
transform 1 0 13156 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_149
timestamp 1636986456
transform 1 0 14260 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 18001
transform 1 0 15364 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 18001
transform 1 0 15916 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1636986456
transform 1 0 16100 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_181
timestamp 1636986456
transform 1 0 17204 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_193
timestamp 1636986456
transform 1 0 18308 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_205
timestamp 1636986456
transform 1 0 19412 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 18001
transform 1 0 20516 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 18001
transform 1 0 21068 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_225
timestamp 1636986456
transform 1 0 21252 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_237
timestamp 1636986456
transform 1 0 22356 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_249
timestamp 1636986456
transform 1 0 23460 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_261
timestamp 1636986456
transform 1 0 24564 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 18001
transform 1 0 25668 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 18001
transform 1 0 26220 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1636986456
transform 1 0 26404 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_293
timestamp 1636986456
transform 1 0 27508 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_305
timestamp 1636986456
transform 1 0 28612 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_317
timestamp 1636986456
transform 1 0 29716 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_329
timestamp 18001
transform 1 0 30820 0 -1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1636986456
transform 1 0 828 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1636986456
transform 1 0 1932 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 18001
transform 1 0 3036 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1636986456
transform 1 0 3220 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1636986456
transform 1 0 4324 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1636986456
transform 1 0 5428 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1636986456
transform 1 0 6532 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 18001
transform 1 0 7636 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 18001
transform 1 0 8188 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1636986456
transform 1 0 8372 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1636986456
transform 1 0 9476 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1636986456
transform 1 0 10580 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1636986456
transform 1 0 11684 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 18001
transform 1 0 12788 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 18001
transform 1 0 13340 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1636986456
transform 1 0 13524 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1636986456
transform 1 0 14628 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_165
timestamp 1636986456
transform 1 0 15732 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_177
timestamp 1636986456
transform 1 0 16836 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 18001
transform 1 0 17940 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 18001
transform 1 0 18492 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1636986456
transform 1 0 18676 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_209
timestamp 1636986456
transform 1 0 19780 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_221
timestamp 1636986456
transform 1 0 20884 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_233
timestamp 1636986456
transform 1 0 21988 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 18001
transform 1 0 23092 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 18001
transform 1 0 23644 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_253
timestamp 1636986456
transform 1 0 23828 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_265
timestamp 1636986456
transform 1 0 24932 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_277
timestamp 1636986456
transform 1 0 26036 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_289
timestamp 1636986456
transform 1 0 27140 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 18001
transform 1 0 28244 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 18001
transform 1 0 28796 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_309
timestamp 1636986456
transform 1 0 28980 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_321
timestamp 18001
transform 1 0 30084 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_329
timestamp 18001
transform 1 0 30820 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1636986456
transform 1 0 828 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1636986456
transform 1 0 1932 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1636986456
transform 1 0 3036 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1636986456
transform 1 0 4140 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 18001
transform 1 0 5244 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 18001
transform 1 0 5612 0 -1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1636986456
transform 1 0 5796 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1636986456
transform 1 0 6900 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1636986456
transform 1 0 8004 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1636986456
transform 1 0 9108 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 18001
transform 1 0 10212 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 18001
transform 1 0 10764 0 -1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1636986456
transform 1 0 10948 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1636986456
transform 1 0 12052 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_137
timestamp 1636986456
transform 1 0 13156 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_149
timestamp 1636986456
transform 1 0 14260 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 18001
transform 1 0 15364 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 18001
transform 1 0 15916 0 -1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1636986456
transform 1 0 16100 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_181
timestamp 1636986456
transform 1 0 17204 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_193
timestamp 1636986456
transform 1 0 18308 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_205
timestamp 1636986456
transform 1 0 19412 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 18001
transform 1 0 20516 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 18001
transform 1 0 21068 0 -1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_225
timestamp 1636986456
transform 1 0 21252 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_237
timestamp 1636986456
transform 1 0 22356 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_249
timestamp 1636986456
transform 1 0 23460 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_261
timestamp 1636986456
transform 1 0 24564 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 18001
transform 1 0 25668 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 18001
transform 1 0 26220 0 -1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_281
timestamp 1636986456
transform 1 0 26404 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_293
timestamp 1636986456
transform 1 0 27508 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_305
timestamp 1636986456
transform 1 0 28612 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_317
timestamp 1636986456
transform 1 0 29716 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_329
timestamp 18001
transform 1 0 30820 0 -1 8160
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1636986456
transform 1 0 828 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1636986456
transform 1 0 1932 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 18001
transform 1 0 3036 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1636986456
transform 1 0 3220 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1636986456
transform 1 0 4324 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1636986456
transform 1 0 5428 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1636986456
transform 1 0 6532 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 18001
transform 1 0 7636 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 18001
transform 1 0 8188 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1636986456
transform 1 0 8372 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1636986456
transform 1 0 9476 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1636986456
transform 1 0 10580 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_121
timestamp 1636986456
transform 1 0 11684 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 18001
transform 1 0 12788 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 18001
transform 1 0 13340 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1636986456
transform 1 0 13524 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1636986456
transform 1 0 14628 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_165
timestamp 1636986456
transform 1 0 15732 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_177
timestamp 1636986456
transform 1 0 16836 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 18001
transform 1 0 17940 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 18001
transform 1 0 18492 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_197
timestamp 1636986456
transform 1 0 18676 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_209
timestamp 1636986456
transform 1 0 19780 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_221
timestamp 1636986456
transform 1 0 20884 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_233
timestamp 1636986456
transform 1 0 21988 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 18001
transform 1 0 23092 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 18001
transform 1 0 23644 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_253
timestamp 1636986456
transform 1 0 23828 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_265
timestamp 1636986456
transform 1 0 24932 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_277
timestamp 1636986456
transform 1 0 26036 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_289
timestamp 1636986456
transform 1 0 27140 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_301
timestamp 18001
transform 1 0 28244 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 18001
transform 1 0 28796 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_309
timestamp 1636986456
transform 1 0 28980 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_321
timestamp 18001
transform 1 0 30084 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_329
timestamp 18001
transform 1 0 30820 0 1 8160
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1636986456
transform 1 0 828 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1636986456
transform 1 0 1932 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1636986456
transform 1 0 3036 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1636986456
transform 1 0 4140 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 18001
transform 1 0 5244 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 18001
transform 1 0 5612 0 -1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1636986456
transform 1 0 5796 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1636986456
transform 1 0 6900 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1636986456
transform 1 0 8004 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1636986456
transform 1 0 9108 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 18001
transform 1 0 10212 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 18001
transform 1 0 10764 0 -1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1636986456
transform 1 0 10948 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_125
timestamp 1636986456
transform 1 0 12052 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_137
timestamp 1636986456
transform 1 0 13156 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_149
timestamp 1636986456
transform 1 0 14260 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 18001
transform 1 0 15364 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 18001
transform 1 0 15916 0 -1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1636986456
transform 1 0 16100 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_181
timestamp 1636986456
transform 1 0 17204 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_193
timestamp 1636986456
transform 1 0 18308 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_205
timestamp 1636986456
transform 1 0 19412 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 18001
transform 1 0 20516 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 18001
transform 1 0 21068 0 -1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_225
timestamp 1636986456
transform 1 0 21252 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_237
timestamp 1636986456
transform 1 0 22356 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_249
timestamp 1636986456
transform 1 0 23460 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_261
timestamp 1636986456
transform 1 0 24564 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_273
timestamp 18001
transform 1 0 25668 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 18001
transform 1 0 26220 0 -1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_281
timestamp 1636986456
transform 1 0 26404 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_293
timestamp 1636986456
transform 1 0 27508 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_305
timestamp 1636986456
transform 1 0 28612 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_317
timestamp 1636986456
transform 1 0 29716 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_329
timestamp 18001
transform 1 0 30820 0 -1 9248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1636986456
transform 1 0 828 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1636986456
transform 1 0 1932 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 18001
transform 1 0 3036 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1636986456
transform 1 0 3220 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1636986456
transform 1 0 4324 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1636986456
transform 1 0 5428 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1636986456
transform 1 0 6532 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 18001
transform 1 0 7636 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 18001
transform 1 0 8188 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1636986456
transform 1 0 8372 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1636986456
transform 1 0 9476 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 1636986456
transform 1 0 10580 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_121
timestamp 1636986456
transform 1 0 11684 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 18001
transform 1 0 12788 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 18001
transform 1 0 13340 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1636986456
transform 1 0 13524 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_153
timestamp 1636986456
transform 1 0 14628 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_165
timestamp 1636986456
transform 1 0 15732 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_177
timestamp 1636986456
transform 1 0 16836 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 18001
transform 1 0 17940 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 18001
transform 1 0 18492 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_197
timestamp 1636986456
transform 1 0 18676 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_209
timestamp 1636986456
transform 1 0 19780 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_221
timestamp 1636986456
transform 1 0 20884 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_233
timestamp 1636986456
transform 1 0 21988 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_245
timestamp 18001
transform 1 0 23092 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 18001
transform 1 0 23644 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_253
timestamp 1636986456
transform 1 0 23828 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_265
timestamp 1636986456
transform 1 0 24932 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_277
timestamp 1636986456
transform 1 0 26036 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_289
timestamp 1636986456
transform 1 0 27140 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_301
timestamp 18001
transform 1 0 28244 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 18001
transform 1 0 28796 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_309
timestamp 1636986456
transform 1 0 28980 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_321
timestamp 18001
transform 1 0 30084 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_329
timestamp 18001
transform 1 0 30820 0 1 9248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1636986456
transform 1 0 828 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1636986456
transform 1 0 1932 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1636986456
transform 1 0 3036 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_39
timestamp 1636986456
transform 1 0 4140 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 18001
transform 1 0 5244 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 18001
transform 1 0 5612 0 -1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1636986456
transform 1 0 5796 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1636986456
transform 1 0 6900 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1636986456
transform 1 0 8004 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1636986456
transform 1 0 9108 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 18001
transform 1 0 10212 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 18001
transform 1 0 10764 0 -1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1636986456
transform 1 0 10948 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_125
timestamp 1636986456
transform 1 0 12052 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_137
timestamp 1636986456
transform 1 0 13156 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_149
timestamp 1636986456
transform 1 0 14260 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 18001
transform 1 0 15364 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 18001
transform 1 0 15916 0 -1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_169
timestamp 1636986456
transform 1 0 16100 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_181
timestamp 1636986456
transform 1 0 17204 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_193
timestamp 1636986456
transform 1 0 18308 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_205
timestamp 1636986456
transform 1 0 19412 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_217
timestamp 18001
transform 1 0 20516 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 18001
transform 1 0 21068 0 -1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_225
timestamp 1636986456
transform 1 0 21252 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_237
timestamp 1636986456
transform 1 0 22356 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_249
timestamp 1636986456
transform 1 0 23460 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_261
timestamp 1636986456
transform 1 0 24564 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 18001
transform 1 0 25668 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 18001
transform 1 0 26220 0 -1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_281
timestamp 1636986456
transform 1 0 26404 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_293
timestamp 1636986456
transform 1 0 27508 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_305
timestamp 1636986456
transform 1 0 28612 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_317
timestamp 1636986456
transform 1 0 29716 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_329
timestamp 18001
transform 1 0 30820 0 -1 10336
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1636986456
transform 1 0 828 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1636986456
transform 1 0 1932 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 18001
transform 1 0 3036 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1636986456
transform 1 0 3220 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1636986456
transform 1 0 4324 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1636986456
transform 1 0 5428 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1636986456
transform 1 0 6532 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 18001
transform 1 0 7636 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 18001
transform 1 0 8188 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1636986456
transform 1 0 8372 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1636986456
transform 1 0 9476 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1636986456
transform 1 0 10580 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_121
timestamp 1636986456
transform 1 0 11684 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 18001
transform 1 0 12788 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 18001
transform 1 0 13340 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1636986456
transform 1 0 13524 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_153
timestamp 1636986456
transform 1 0 14628 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_165
timestamp 1636986456
transform 1 0 15732 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_177
timestamp 1636986456
transform 1 0 16836 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 18001
transform 1 0 17940 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 18001
transform 1 0 18492 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_197
timestamp 1636986456
transform 1 0 18676 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_209
timestamp 1636986456
transform 1 0 19780 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_221
timestamp 1636986456
transform 1 0 20884 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_233
timestamp 1636986456
transform 1 0 21988 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_245
timestamp 18001
transform 1 0 23092 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 18001
transform 1 0 23644 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_253
timestamp 1636986456
transform 1 0 23828 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_265
timestamp 1636986456
transform 1 0 24932 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_277
timestamp 1636986456
transform 1 0 26036 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_289
timestamp 1636986456
transform 1 0 27140 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_301
timestamp 18001
transform 1 0 28244 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 18001
transform 1 0 28796 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_309
timestamp 1636986456
transform 1 0 28980 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_321
timestamp 18001
transform 1 0 30084 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_329
timestamp 18001
transform 1 0 30820 0 1 10336
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1636986456
transform 1 0 828 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1636986456
transform 1 0 1932 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1636986456
transform 1 0 3036 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1636986456
transform 1 0 4140 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 18001
transform 1 0 5244 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 18001
transform 1 0 5612 0 -1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1636986456
transform 1 0 5796 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1636986456
transform 1 0 6900 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1636986456
transform 1 0 8004 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1636986456
transform 1 0 9108 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 18001
transform 1 0 10212 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 18001
transform 1 0 10764 0 -1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1636986456
transform 1 0 10948 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_125
timestamp 1636986456
transform 1 0 12052 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_137
timestamp 1636986456
transform 1 0 13156 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_149
timestamp 1636986456
transform 1 0 14260 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 18001
transform 1 0 15364 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 18001
transform 1 0 15916 0 -1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_169
timestamp 1636986456
transform 1 0 16100 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_181
timestamp 1636986456
transform 1 0 17204 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_193
timestamp 1636986456
transform 1 0 18308 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_205
timestamp 1636986456
transform 1 0 19412 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_217
timestamp 18001
transform 1 0 20516 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 18001
transform 1 0 21068 0 -1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_225
timestamp 1636986456
transform 1 0 21252 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_237
timestamp 1636986456
transform 1 0 22356 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_249
timestamp 1636986456
transform 1 0 23460 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_261
timestamp 1636986456
transform 1 0 24564 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_273
timestamp 18001
transform 1 0 25668 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 18001
transform 1 0 26220 0 -1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_281
timestamp 1636986456
transform 1 0 26404 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_293
timestamp 1636986456
transform 1 0 27508 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_305
timestamp 1636986456
transform 1 0 28612 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_317
timestamp 1636986456
transform 1 0 29716 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_329
timestamp 18001
transform 1 0 30820 0 -1 11424
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1636986456
transform 1 0 828 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1636986456
transform 1 0 1932 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 18001
transform 1 0 3036 0 1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1636986456
transform 1 0 3220 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1636986456
transform 1 0 4324 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1636986456
transform 1 0 5428 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1636986456
transform 1 0 6532 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 18001
transform 1 0 7636 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 18001
transform 1 0 8188 0 1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1636986456
transform 1 0 8372 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_97
timestamp 1636986456
transform 1 0 9476 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_109
timestamp 1636986456
transform 1 0 10580 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_121
timestamp 1636986456
transform 1 0 11684 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 18001
transform 1 0 12788 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 18001
transform 1 0 13340 0 1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1636986456
transform 1 0 13524 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_153
timestamp 1636986456
transform 1 0 14628 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_165
timestamp 1636986456
transform 1 0 15732 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_177
timestamp 1636986456
transform 1 0 16836 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_189
timestamp 18001
transform 1 0 17940 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 18001
transform 1 0 18492 0 1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_197
timestamp 1636986456
transform 1 0 18676 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_209
timestamp 1636986456
transform 1 0 19780 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_221
timestamp 1636986456
transform 1 0 20884 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_233
timestamp 1636986456
transform 1 0 21988 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_245
timestamp 18001
transform 1 0 23092 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 18001
transform 1 0 23644 0 1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_253
timestamp 1636986456
transform 1 0 23828 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_265
timestamp 1636986456
transform 1 0 24932 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_277
timestamp 1636986456
transform 1 0 26036 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_289
timestamp 1636986456
transform 1 0 27140 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_301
timestamp 18001
transform 1 0 28244 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 18001
transform 1 0 28796 0 1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_309
timestamp 1636986456
transform 1 0 28980 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_321
timestamp 18001
transform 1 0 30084 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_329
timestamp 18001
transform 1 0 30820 0 1 11424
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1636986456
transform 1 0 828 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1636986456
transform 1 0 1932 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_27
timestamp 1636986456
transform 1 0 3036 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_39
timestamp 1636986456
transform 1 0 4140 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 18001
transform 1 0 5244 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 18001
transform 1 0 5612 0 -1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1636986456
transform 1 0 5796 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1636986456
transform 1 0 6900 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_81
timestamp 1636986456
transform 1 0 8004 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_93
timestamp 1636986456
transform 1 0 9108 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 18001
transform 1 0 10212 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 18001
transform 1 0 10764 0 -1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1636986456
transform 1 0 10948 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_125
timestamp 1636986456
transform 1 0 12052 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_137
timestamp 1636986456
transform 1 0 13156 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_149
timestamp 1636986456
transform 1 0 14260 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 18001
transform 1 0 15364 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 18001
transform 1 0 15916 0 -1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_169
timestamp 1636986456
transform 1 0 16100 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_181
timestamp 1636986456
transform 1 0 17204 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_193
timestamp 1636986456
transform 1 0 18308 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_205
timestamp 1636986456
transform 1 0 19412 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_217
timestamp 18001
transform 1 0 20516 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 18001
transform 1 0 21068 0 -1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_225
timestamp 1636986456
transform 1 0 21252 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_237
timestamp 1636986456
transform 1 0 22356 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_249
timestamp 1636986456
transform 1 0 23460 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_261
timestamp 1636986456
transform 1 0 24564 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_273
timestamp 18001
transform 1 0 25668 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 18001
transform 1 0 26220 0 -1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_281
timestamp 1636986456
transform 1 0 26404 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_293
timestamp 1636986456
transform 1 0 27508 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_305
timestamp 1636986456
transform 1 0 28612 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_317
timestamp 1636986456
transform 1 0 29716 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_329
timestamp 18001
transform 1 0 30820 0 -1 12512
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1636986456
transform 1 0 828 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1636986456
transform 1 0 1932 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 18001
transform 1 0 3036 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1636986456
transform 1 0 3220 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1636986456
transform 1 0 4324 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1636986456
transform 1 0 5428 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1636986456
transform 1 0 6532 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 18001
transform 1 0 7636 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 18001
transform 1 0 8188 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1636986456
transform 1 0 8372 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_97
timestamp 1636986456
transform 1 0 9476 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_109
timestamp 1636986456
transform 1 0 10580 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_121
timestamp 1636986456
transform 1 0 11684 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 18001
transform 1 0 12788 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 18001
transform 1 0 13340 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1636986456
transform 1 0 13524 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_153
timestamp 1636986456
transform 1 0 14628 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_165
timestamp 1636986456
transform 1 0 15732 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_177
timestamp 1636986456
transform 1 0 16836 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_189
timestamp 18001
transform 1 0 17940 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 18001
transform 1 0 18492 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_197
timestamp 1636986456
transform 1 0 18676 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_209
timestamp 1636986456
transform 1 0 19780 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_221
timestamp 1636986456
transform 1 0 20884 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_233
timestamp 1636986456
transform 1 0 21988 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_245
timestamp 18001
transform 1 0 23092 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 18001
transform 1 0 23644 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_253
timestamp 1636986456
transform 1 0 23828 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_265
timestamp 1636986456
transform 1 0 24932 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_277
timestamp 1636986456
transform 1 0 26036 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_289
timestamp 1636986456
transform 1 0 27140 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_301
timestamp 18001
transform 1 0 28244 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 18001
transform 1 0 28796 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_309
timestamp 1636986456
transform 1 0 28980 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_321
timestamp 18001
transform 1 0 30084 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_329
timestamp 18001
transform 1 0 30820 0 1 12512
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1636986456
transform 1 0 828 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1636986456
transform 1 0 1932 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1636986456
transform 1 0 3036 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1636986456
transform 1 0 4140 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 18001
transform 1 0 5244 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 18001
transform 1 0 5612 0 -1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1636986456
transform 1 0 5796 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1636986456
transform 1 0 6900 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_81
timestamp 1636986456
transform 1 0 8004 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_93
timestamp 1636986456
transform 1 0 9108 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 18001
transform 1 0 10212 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 18001
transform 1 0 10764 0 -1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1636986456
transform 1 0 10948 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_125
timestamp 1636986456
transform 1 0 12052 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_137
timestamp 1636986456
transform 1 0 13156 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_149
timestamp 1636986456
transform 1 0 14260 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 18001
transform 1 0 15364 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 18001
transform 1 0 15916 0 -1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_169
timestamp 1636986456
transform 1 0 16100 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_181
timestamp 1636986456
transform 1 0 17204 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_193
timestamp 1636986456
transform 1 0 18308 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_205
timestamp 1636986456
transform 1 0 19412 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_217
timestamp 18001
transform 1 0 20516 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 18001
transform 1 0 21068 0 -1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_225
timestamp 1636986456
transform 1 0 21252 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_237
timestamp 1636986456
transform 1 0 22356 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_249
timestamp 1636986456
transform 1 0 23460 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_261
timestamp 1636986456
transform 1 0 24564 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_273
timestamp 18001
transform 1 0 25668 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 18001
transform 1 0 26220 0 -1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_281
timestamp 1636986456
transform 1 0 26404 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_293
timestamp 1636986456
transform 1 0 27508 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_305
timestamp 1636986456
transform 1 0 28612 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_317
timestamp 1636986456
transform 1 0 29716 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_329
timestamp 18001
transform 1 0 30820 0 -1 13600
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1636986456
transform 1 0 828 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1636986456
transform 1 0 1932 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 18001
transform 1 0 3036 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1636986456
transform 1 0 3220 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1636986456
transform 1 0 4324 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1636986456
transform 1 0 5428 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1636986456
transform 1 0 6532 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 18001
transform 1 0 7636 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 18001
transform 1 0 8188 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1636986456
transform 1 0 8372 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_97
timestamp 1636986456
transform 1 0 9476 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_109
timestamp 1636986456
transform 1 0 10580 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_121
timestamp 1636986456
transform 1 0 11684 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 18001
transform 1 0 12788 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 18001
transform 1 0 13340 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_161
timestamp 1636986456
transform 1 0 15364 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_173
timestamp 18001
transform 1 0 16468 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_186
timestamp 18001
transform 1 0 17664 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_194
timestamp 18001
transform 1 0 18400 0 1 13600
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_197
timestamp 1636986456
transform 1 0 18676 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_209
timestamp 1636986456
transform 1 0 19780 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_221
timestamp 1636986456
transform 1 0 20884 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_233
timestamp 1636986456
transform 1 0 21988 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_245
timestamp 18001
transform 1 0 23092 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 18001
transform 1 0 23644 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_253
timestamp 1636986456
transform 1 0 23828 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_265
timestamp 1636986456
transform 1 0 24932 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_277
timestamp 1636986456
transform 1 0 26036 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_289
timestamp 1636986456
transform 1 0 27140 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_301
timestamp 18001
transform 1 0 28244 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 18001
transform 1 0 28796 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_309
timestamp 1636986456
transform 1 0 28980 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_321
timestamp 18001
transform 1 0 30084 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_329
timestamp 18001
transform 1 0 30820 0 1 13600
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1636986456
transform 1 0 828 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1636986456
transform 1 0 1932 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_27
timestamp 1636986456
transform 1 0 3036 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_39
timestamp 1636986456
transform 1 0 4140 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 18001
transform 1 0 5244 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 18001
transform 1 0 5612 0 -1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1636986456
transform 1 0 5796 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1636986456
transform 1 0 6900 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_81
timestamp 1636986456
transform 1 0 8004 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_93
timestamp 1636986456
transform 1 0 9108 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 18001
transform 1 0 10212 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 18001
transform 1 0 10764 0 -1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1636986456
transform 1 0 10948 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_125
timestamp 18001
transform 1 0 12052 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_131
timestamp 18001
transform 1 0 12604 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_157
timestamp 18001
transform 1 0 14996 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_165
timestamp 18001
transform 1 0 15732 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_169
timestamp 18001
transform 1 0 16100 0 -1 14688
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_199
timestamp 1636986456
transform 1 0 18860 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_211
timestamp 1636986456
transform 1 0 19964 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 18001
transform 1 0 21068 0 -1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_225
timestamp 1636986456
transform 1 0 21252 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_237
timestamp 1636986456
transform 1 0 22356 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_249
timestamp 1636986456
transform 1 0 23460 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_261
timestamp 1636986456
transform 1 0 24564 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_273
timestamp 18001
transform 1 0 25668 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 18001
transform 1 0 26220 0 -1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_281
timestamp 1636986456
transform 1 0 26404 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_293
timestamp 1636986456
transform 1 0 27508 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_305
timestamp 1636986456
transform 1 0 28612 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_317
timestamp 1636986456
transform 1 0 29716 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1636986456
transform 1 0 828 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1636986456
transform 1 0 1932 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 18001
transform 1 0 3036 0 1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1636986456
transform 1 0 3220 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1636986456
transform 1 0 4324 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1636986456
transform 1 0 5428 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_65
timestamp 1636986456
transform 1 0 6532 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 18001
transform 1 0 7636 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 18001
transform 1 0 8188 0 1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1636986456
transform 1 0 8372 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 1636986456
transform 1 0 9476 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_109
timestamp 1636986456
transform 1 0 10580 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_121
timestamp 18001
transform 1 0 11684 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_127
timestamp 18001
transform 1 0 12236 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_146
timestamp 18001
transform 1 0 13984 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_168
timestamp 18001
transform 1 0 16008 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_26_187
timestamp 18001
transform 1 0 17756 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 18001
transform 1 0 18492 0 1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_197
timestamp 1636986456
transform 1 0 18676 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_209
timestamp 1636986456
transform 1 0 19780 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_221
timestamp 1636986456
transform 1 0 20884 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_233
timestamp 1636986456
transform 1 0 21988 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_245
timestamp 18001
transform 1 0 23092 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 18001
transform 1 0 23644 0 1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_253
timestamp 1636986456
transform 1 0 23828 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_265
timestamp 1636986456
transform 1 0 24932 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_277
timestamp 1636986456
transform 1 0 26036 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_289
timestamp 1636986456
transform 1 0 27140 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_301
timestamp 18001
transform 1 0 28244 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 18001
transform 1 0 28796 0 1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_309
timestamp 1636986456
transform 1 0 28980 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_321
timestamp 18001
transform 1 0 30084 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_329
timestamp 18001
transform 1 0 30820 0 1 14688
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1636986456
transform 1 0 828 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1636986456
transform 1 0 1932 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_27
timestamp 1636986456
transform 1 0 3036 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_39
timestamp 1636986456
transform 1 0 4140 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 18001
transform 1 0 5244 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 18001
transform 1 0 5612 0 -1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1636986456
transform 1 0 5796 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1636986456
transform 1 0 6900 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_81
timestamp 1636986456
transform 1 0 8004 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_93
timestamp 1636986456
transform 1 0 9108 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 18001
transform 1 0 10212 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 18001
transform 1 0 10764 0 -1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1636986456
transform 1 0 10948 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_125
timestamp 18001
transform 1 0 12052 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_160
timestamp 18001
transform 1 0 15272 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_164
timestamp 18001
transform 1 0 15640 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_169
timestamp 18001
transform 1 0 16100 0 -1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_205
timestamp 1636986456
transform 1 0 19412 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_217
timestamp 18001
transform 1 0 20516 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 18001
transform 1 0 21068 0 -1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_225
timestamp 1636986456
transform 1 0 21252 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_237
timestamp 1636986456
transform 1 0 22356 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_249
timestamp 1636986456
transform 1 0 23460 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_261
timestamp 1636986456
transform 1 0 24564 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_273
timestamp 18001
transform 1 0 25668 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 18001
transform 1 0 26220 0 -1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_281
timestamp 1636986456
transform 1 0 26404 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_293
timestamp 1636986456
transform 1 0 27508 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_305
timestamp 1636986456
transform 1 0 28612 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_317
timestamp 1636986456
transform 1 0 29716 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_329
timestamp 18001
transform 1 0 30820 0 -1 15776
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1636986456
transform 1 0 828 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1636986456
transform 1 0 1932 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 18001
transform 1 0 3036 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1636986456
transform 1 0 3220 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1636986456
transform 1 0 4324 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1636986456
transform 1 0 5428 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_65
timestamp 1636986456
transform 1 0 6532 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 18001
transform 1 0 7636 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 18001
transform 1 0 8188 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1636986456
transform 1 0 8372 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_97
timestamp 1636986456
transform 1 0 9476 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_109
timestamp 1636986456
transform 1 0 10580 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_121
timestamp 18001
transform 1 0 11684 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_129
timestamp 18001
transform 1 0 12420 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 18001
transform 1 0 13340 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_148
timestamp 18001
transform 1 0 14168 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_156
timestamp 18001
transform 1 0 14904 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_197
timestamp 1636986456
transform 1 0 18676 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_209
timestamp 1636986456
transform 1 0 19780 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_221
timestamp 1636986456
transform 1 0 20884 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_233
timestamp 1636986456
transform 1 0 21988 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_245
timestamp 18001
transform 1 0 23092 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 18001
transform 1 0 23644 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_253
timestamp 1636986456
transform 1 0 23828 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_265
timestamp 1636986456
transform 1 0 24932 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_277
timestamp 1636986456
transform 1 0 26036 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_289
timestamp 1636986456
transform 1 0 27140 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_301
timestamp 18001
transform 1 0 28244 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp 18001
transform 1 0 28796 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_309
timestamp 1636986456
transform 1 0 28980 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_321
timestamp 18001
transform 1 0 30084 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_329
timestamp 18001
transform 1 0 30820 0 1 15776
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1636986456
transform 1 0 828 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_15
timestamp 1636986456
transform 1 0 1932 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_27
timestamp 1636986456
transform 1 0 3036 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_39
timestamp 1636986456
transform 1 0 4140 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 18001
transform 1 0 5244 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 18001
transform 1 0 5612 0 -1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1636986456
transform 1 0 5796 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_69
timestamp 1636986456
transform 1 0 6900 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_81
timestamp 1636986456
transform 1 0 8004 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_93
timestamp 1636986456
transform 1 0 9108 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 18001
transform 1 0 10212 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 18001
transform 1 0 10764 0 -1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 1636986456
transform 1 0 10948 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_125
timestamp 18001
transform 1 0 12052 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_131
timestamp 18001
transform 1 0 12604 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_164
timestamp 18001
transform 1 0 15640 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_182
timestamp 18001
transform 1 0 17296 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 18001
transform 1 0 21068 0 -1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_225
timestamp 1636986456
transform 1 0 21252 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_237
timestamp 1636986456
transform 1 0 22356 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_249
timestamp 1636986456
transform 1 0 23460 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_261
timestamp 1636986456
transform 1 0 24564 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_273
timestamp 18001
transform 1 0 25668 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp 18001
transform 1 0 26220 0 -1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_281
timestamp 1636986456
transform 1 0 26404 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_293
timestamp 1636986456
transform 1 0 27508 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_305
timestamp 1636986456
transform 1 0 28612 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_317
timestamp 1636986456
transform 1 0 29716 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_329
timestamp 18001
transform 1 0 30820 0 -1 16864
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1636986456
transform 1 0 828 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1636986456
transform 1 0 1932 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 18001
transform 1 0 3036 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1636986456
transform 1 0 3220 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1636986456
transform 1 0 4324 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1636986456
transform 1 0 5428 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_65
timestamp 1636986456
transform 1 0 6532 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 18001
transform 1 0 7636 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 18001
transform 1 0 8188 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1636986456
transform 1 0 8372 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_97
timestamp 1636986456
transform 1 0 9476 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_109
timestamp 1636986456
transform 1 0 10580 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_121
timestamp 18001
transform 1 0 11684 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_129
timestamp 18001
transform 1 0 12420 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_138
timestamp 18001
transform 1 0 13248 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_141
timestamp 18001
transform 1 0 13524 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_149
timestamp 18001
transform 1 0 14260 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_153
timestamp 18001
transform 1 0 14628 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_197
timestamp 1636986456
transform 1 0 18676 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_209
timestamp 1636986456
transform 1 0 19780 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_221
timestamp 1636986456
transform 1 0 20884 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_233
timestamp 1636986456
transform 1 0 21988 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_245
timestamp 18001
transform 1 0 23092 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_251
timestamp 18001
transform 1 0 23644 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_253
timestamp 1636986456
transform 1 0 23828 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_265
timestamp 1636986456
transform 1 0 24932 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_277
timestamp 1636986456
transform 1 0 26036 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_289
timestamp 1636986456
transform 1 0 27140 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_301
timestamp 18001
transform 1 0 28244 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_307
timestamp 18001
transform 1 0 28796 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_309
timestamp 1636986456
transform 1 0 28980 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_321
timestamp 18001
transform 1 0 30084 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_329
timestamp 18001
transform 1 0 30820 0 1 16864
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1636986456
transform 1 0 828 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1636986456
transform 1 0 1932 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_27
timestamp 1636986456
transform 1 0 3036 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_39
timestamp 1636986456
transform 1 0 4140 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 18001
transform 1 0 5244 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 18001
transform 1 0 5612 0 -1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1636986456
transform 1 0 5796 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 1636986456
transform 1 0 6900 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_81
timestamp 1636986456
transform 1 0 8004 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_93
timestamp 1636986456
transform 1 0 9108 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 18001
transform 1 0 10212 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 18001
transform 1 0 10764 0 -1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_113
timestamp 1636986456
transform 1 0 10948 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_125
timestamp 18001
transform 1 0 12052 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_152
timestamp 18001
transform 1 0 14536 0 -1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_204
timestamp 1636986456
transform 1 0 19320 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_216
timestamp 18001
transform 1 0 20424 0 -1 17952
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_31_225
timestamp 1636986456
transform 1 0 21252 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_237
timestamp 1636986456
transform 1 0 22356 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_249
timestamp 1636986456
transform 1 0 23460 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_261
timestamp 1636986456
transform 1 0 24564 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_273
timestamp 18001
transform 1 0 25668 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 18001
transform 1 0 26220 0 -1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_281
timestamp 1636986456
transform 1 0 26404 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_293
timestamp 1636986456
transform 1 0 27508 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_305
timestamp 1636986456
transform 1 0 28612 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_317
timestamp 1636986456
transform 1 0 29716 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_329
timestamp 18001
transform 1 0 30820 0 -1 17952
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1636986456
transform 1 0 828 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_15
timestamp 1636986456
transform 1 0 1932 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 18001
transform 1 0 3036 0 1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1636986456
transform 1 0 3220 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1636986456
transform 1 0 4324 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_53
timestamp 1636986456
transform 1 0 5428 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_65
timestamp 1636986456
transform 1 0 6532 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 18001
transform 1 0 7636 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 18001
transform 1 0 8188 0 1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 1636986456
transform 1 0 8372 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_97
timestamp 1636986456
transform 1 0 9476 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_109
timestamp 1636986456
transform 1 0 10580 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_121
timestamp 1636986456
transform 1 0 11684 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_133
timestamp 18001
transform 1 0 12788 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 18001
transform 1 0 13340 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_161
timestamp 18001
transform 1 0 15364 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_192
timestamp 18001
transform 1 0 18216 0 1 17952
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_197
timestamp 1636986456
transform 1 0 18676 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_209
timestamp 1636986456
transform 1 0 19780 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_221
timestamp 1636986456
transform 1 0 20884 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_233
timestamp 1636986456
transform 1 0 21988 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_245
timestamp 18001
transform 1 0 23092 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 18001
transform 1 0 23644 0 1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_253
timestamp 1636986456
transform 1 0 23828 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_265
timestamp 1636986456
transform 1 0 24932 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_277
timestamp 1636986456
transform 1 0 26036 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_289
timestamp 1636986456
transform 1 0 27140 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_301
timestamp 18001
transform 1 0 28244 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_307
timestamp 18001
transform 1 0 28796 0 1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_309
timestamp 1636986456
transform 1 0 28980 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_321
timestamp 18001
transform 1 0 30084 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_329
timestamp 18001
transform 1 0 30820 0 1 17952
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_6
timestamp 1636986456
transform 1 0 1104 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_18
timestamp 18001
transform 1 0 2208 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_26
timestamp 18001
transform 1 0 2944 0 -1 19040
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_29
timestamp 1636986456
transform 1 0 3220 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_41
timestamp 1636986456
transform 1 0 4324 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_53
timestamp 18001
transform 1 0 5428 0 -1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1636986456
transform 1 0 5796 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_69
timestamp 1636986456
transform 1 0 6900 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_81
timestamp 18001
transform 1 0 8004 0 -1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_85
timestamp 1636986456
transform 1 0 8372 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_97
timestamp 18001
transform 1 0 9476 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_105
timestamp 18001
transform 1 0 10212 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_110
timestamp 18001
transform 1 0 10672 0 -1 19040
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1636986456
transform 1 0 10948 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_125
timestamp 18001
transform 1 0 12052 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_131
timestamp 18001
transform 1 0 12604 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_138
timestamp 18001
transform 1 0 13248 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_141
timestamp 18001
transform 1 0 13524 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_145
timestamp 18001
transform 1 0 13892 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_152
timestamp 18001
transform 1 0 14536 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_157
timestamp 18001
transform 1 0 14996 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 18001
transform 1 0 15916 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_177
timestamp 18001
transform 1 0 16836 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_194
timestamp 18001
transform 1 0 18400 0 -1 19040
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_200
timestamp 1636986456
transform 1 0 18952 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_212
timestamp 1636986456
transform 1 0 20056 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_225
timestamp 1636986456
transform 1 0 21252 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_237
timestamp 18001
transform 1 0 22356 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_33_243
timestamp 18001
transform 1 0 22908 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_251
timestamp 18001
transform 1 0 23644 0 -1 19040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_253
timestamp 1636986456
transform 1 0 23828 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_265
timestamp 1636986456
transform 1 0 24932 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_277
timestamp 18001
transform 1 0 26036 0 -1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_281
timestamp 1636986456
transform 1 0 26404 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_293
timestamp 1636986456
transform 1 0 27508 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_305
timestamp 18001
transform 1 0 28612 0 -1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_309
timestamp 1636986456
transform 1 0 28980 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_321
timestamp 18001
transform 1 0 30084 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_329
timestamp 18001
transform 1 0 30820 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1
timestamp 18001
transform -1 0 14904 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 18001
transform -1 0 15916 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 18001
transform -1 0 16008 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 18001
transform -1 0 18124 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 18001
transform 1 0 17020 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 18001
transform -1 0 17572 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 18001
transform -1 0 16836 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  input1
timestamp 18001
transform 1 0 16836 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 18001
transform -1 0 14536 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_34
timestamp 18001
transform 1 0 552 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 18001
transform -1 0 31372 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_35
timestamp 18001
transform 1 0 552 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 18001
transform -1 0 31372 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_36
timestamp 18001
transform 1 0 552 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 18001
transform -1 0 31372 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_37
timestamp 18001
transform 1 0 552 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 18001
transform -1 0 31372 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_38
timestamp 18001
transform 1 0 552 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 18001
transform -1 0 31372 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_39
timestamp 18001
transform 1 0 552 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 18001
transform -1 0 31372 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_40
timestamp 18001
transform 1 0 552 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 18001
transform -1 0 31372 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_41
timestamp 18001
transform 1 0 552 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 18001
transform -1 0 31372 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_42
timestamp 18001
transform 1 0 552 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 18001
transform -1 0 31372 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_43
timestamp 18001
transform 1 0 552 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 18001
transform -1 0 31372 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_44
timestamp 18001
transform 1 0 552 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 18001
transform -1 0 31372 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_45
timestamp 18001
transform 1 0 552 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 18001
transform -1 0 31372 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_46
timestamp 18001
transform 1 0 552 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 18001
transform -1 0 31372 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_47
timestamp 18001
transform 1 0 552 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 18001
transform -1 0 31372 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_48
timestamp 18001
transform 1 0 552 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 18001
transform -1 0 31372 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_49
timestamp 18001
transform 1 0 552 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 18001
transform -1 0 31372 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_50
timestamp 18001
transform 1 0 552 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 18001
transform -1 0 31372 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_51
timestamp 18001
transform 1 0 552 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 18001
transform -1 0 31372 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_52
timestamp 18001
transform 1 0 552 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 18001
transform -1 0 31372 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_53
timestamp 18001
transform 1 0 552 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 18001
transform -1 0 31372 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_54
timestamp 18001
transform 1 0 552 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 18001
transform -1 0 31372 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_55
timestamp 18001
transform 1 0 552 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 18001
transform -1 0 31372 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_56
timestamp 18001
transform 1 0 552 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 18001
transform -1 0 31372 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_57
timestamp 18001
transform 1 0 552 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 18001
transform -1 0 31372 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_58
timestamp 18001
transform 1 0 552 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 18001
transform -1 0 31372 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_59
timestamp 18001
transform 1 0 552 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 18001
transform -1 0 31372 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_60
timestamp 18001
transform 1 0 552 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 18001
transform -1 0 31372 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_61
timestamp 18001
transform 1 0 552 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 18001
transform -1 0 31372 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_62
timestamp 18001
transform 1 0 552 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 18001
transform -1 0 31372 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_63
timestamp 18001
transform 1 0 552 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp 18001
transform -1 0 31372 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_64
timestamp 18001
transform 1 0 552 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp 18001
transform -1 0 31372 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_65
timestamp 18001
transform 1 0 552 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp 18001
transform -1 0 31372 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_66
timestamp 18001
transform 1 0 552 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp 18001
transform -1 0 31372 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Left_67
timestamp 18001
transform 1 0 552 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Right_33
timestamp 18001
transform -1 0 31372 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  stoplight_example_5
timestamp 18001
transform -1 0 17756 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  stoplight_example_6
timestamp 18001
transform -1 0 19044 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  stoplight_example_7
timestamp 18001
transform -1 0 11960 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  stoplight_example_8
timestamp 18001
transform -1 0 12604 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  stoplight_example_9
timestamp 18001
transform -1 0 13892 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  stoplight_example_10
timestamp 18001
transform -1 0 13892 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  stoplight_example_11
timestamp 18001
transform -1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  stoplight_example_12
timestamp 18001
transform -1 0 14536 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  stoplight_example_13
timestamp 18001
transform -1 0 12604 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  stoplight_example_14
timestamp 18001
transform -1 0 20332 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  stoplight_example_15
timestamp 18001
transform -1 0 10672 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  stoplight_example_16
timestamp 18001
transform -1 0 15824 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  stoplight_example_17
timestamp 18001
transform 1 0 30820 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  stoplight_example_18
timestamp 18001
transform -1 0 7452 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  stoplight_example_19
timestamp 18001
transform -1 0 9384 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  stoplight_example_20
timestamp 18001
transform -1 0 18952 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  stoplight_example_21
timestamp 18001
transform -1 0 22908 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  stoplight_example_22
timestamp 18001
transform -1 0 13248 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  stoplight_example_23
timestamp 18001
transform -1 0 18400 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  stoplight_example_24
timestamp 18001
transform -1 0 15180 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  stoplight_example_25
timestamp 18001
transform -1 0 13248 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_68
timestamp 18001
transform 1 0 3128 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_69
timestamp 18001
transform 1 0 5704 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_70
timestamp 18001
transform 1 0 8280 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_71
timestamp 18001
transform 1 0 10856 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_72
timestamp 18001
transform 1 0 13432 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_73
timestamp 18001
transform 1 0 16008 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_74
timestamp 18001
transform 1 0 18584 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_75
timestamp 18001
transform 1 0 21160 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_76
timestamp 18001
transform 1 0 23736 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_77
timestamp 18001
transform 1 0 26312 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_78
timestamp 18001
transform 1 0 28888 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_79
timestamp 18001
transform 1 0 5704 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_80
timestamp 18001
transform 1 0 10856 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_81
timestamp 18001
transform 1 0 16008 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_82
timestamp 18001
transform 1 0 21160 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_83
timestamp 18001
transform 1 0 26312 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_84
timestamp 18001
transform 1 0 3128 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_85
timestamp 18001
transform 1 0 8280 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_86
timestamp 18001
transform 1 0 13432 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_87
timestamp 18001
transform 1 0 18584 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_88
timestamp 18001
transform 1 0 23736 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_89
timestamp 18001
transform 1 0 28888 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_90
timestamp 18001
transform 1 0 5704 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_91
timestamp 18001
transform 1 0 10856 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_92
timestamp 18001
transform 1 0 16008 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_93
timestamp 18001
transform 1 0 21160 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_94
timestamp 18001
transform 1 0 26312 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_95
timestamp 18001
transform 1 0 3128 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_96
timestamp 18001
transform 1 0 8280 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_97
timestamp 18001
transform 1 0 13432 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_98
timestamp 18001
transform 1 0 18584 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_99
timestamp 18001
transform 1 0 23736 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_100
timestamp 18001
transform 1 0 28888 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_101
timestamp 18001
transform 1 0 5704 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_102
timestamp 18001
transform 1 0 10856 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_103
timestamp 18001
transform 1 0 16008 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_104
timestamp 18001
transform 1 0 21160 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_105
timestamp 18001
transform 1 0 26312 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_106
timestamp 18001
transform 1 0 3128 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_107
timestamp 18001
transform 1 0 8280 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_108
timestamp 18001
transform 1 0 13432 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_109
timestamp 18001
transform 1 0 18584 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_110
timestamp 18001
transform 1 0 23736 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_111
timestamp 18001
transform 1 0 28888 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_112
timestamp 18001
transform 1 0 5704 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_113
timestamp 18001
transform 1 0 10856 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_114
timestamp 18001
transform 1 0 16008 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_115
timestamp 18001
transform 1 0 21160 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_116
timestamp 18001
transform 1 0 26312 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_117
timestamp 18001
transform 1 0 3128 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_118
timestamp 18001
transform 1 0 8280 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_119
timestamp 18001
transform 1 0 13432 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_120
timestamp 18001
transform 1 0 18584 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_121
timestamp 18001
transform 1 0 23736 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_122
timestamp 18001
transform 1 0 28888 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_123
timestamp 18001
transform 1 0 5704 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_124
timestamp 18001
transform 1 0 10856 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_125
timestamp 18001
transform 1 0 16008 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_126
timestamp 18001
transform 1 0 21160 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_127
timestamp 18001
transform 1 0 26312 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_128
timestamp 18001
transform 1 0 3128 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_129
timestamp 18001
transform 1 0 8280 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_130
timestamp 18001
transform 1 0 13432 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_131
timestamp 18001
transform 1 0 18584 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_132
timestamp 18001
transform 1 0 23736 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_133
timestamp 18001
transform 1 0 28888 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_134
timestamp 18001
transform 1 0 5704 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_135
timestamp 18001
transform 1 0 10856 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_136
timestamp 18001
transform 1 0 16008 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_137
timestamp 18001
transform 1 0 21160 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_138
timestamp 18001
transform 1 0 26312 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_139
timestamp 18001
transform 1 0 3128 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_140
timestamp 18001
transform 1 0 8280 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_141
timestamp 18001
transform 1 0 13432 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_142
timestamp 18001
transform 1 0 18584 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_143
timestamp 18001
transform 1 0 23736 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_144
timestamp 18001
transform 1 0 28888 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_145
timestamp 18001
transform 1 0 5704 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_146
timestamp 18001
transform 1 0 10856 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_147
timestamp 18001
transform 1 0 16008 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_148
timestamp 18001
transform 1 0 21160 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_149
timestamp 18001
transform 1 0 26312 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_150
timestamp 18001
transform 1 0 3128 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_151
timestamp 18001
transform 1 0 8280 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_152
timestamp 18001
transform 1 0 13432 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_153
timestamp 18001
transform 1 0 18584 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_154
timestamp 18001
transform 1 0 23736 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_155
timestamp 18001
transform 1 0 28888 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_156
timestamp 18001
transform 1 0 5704 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_157
timestamp 18001
transform 1 0 10856 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_158
timestamp 18001
transform 1 0 16008 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_159
timestamp 18001
transform 1 0 21160 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_160
timestamp 18001
transform 1 0 26312 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_161
timestamp 18001
transform 1 0 3128 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_162
timestamp 18001
transform 1 0 8280 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_163
timestamp 18001
transform 1 0 13432 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_164
timestamp 18001
transform 1 0 18584 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_165
timestamp 18001
transform 1 0 23736 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_166
timestamp 18001
transform 1 0 28888 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_167
timestamp 18001
transform 1 0 5704 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_168
timestamp 18001
transform 1 0 10856 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_169
timestamp 18001
transform 1 0 16008 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_170
timestamp 18001
transform 1 0 21160 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_171
timestamp 18001
transform 1 0 26312 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_172
timestamp 18001
transform 1 0 3128 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_173
timestamp 18001
transform 1 0 8280 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_174
timestamp 18001
transform 1 0 13432 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_175
timestamp 18001
transform 1 0 18584 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_176
timestamp 18001
transform 1 0 23736 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_177
timestamp 18001
transform 1 0 28888 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_178
timestamp 18001
transform 1 0 5704 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_179
timestamp 18001
transform 1 0 10856 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_180
timestamp 18001
transform 1 0 16008 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_181
timestamp 18001
transform 1 0 21160 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_182
timestamp 18001
transform 1 0 26312 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_183
timestamp 18001
transform 1 0 3128 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_184
timestamp 18001
transform 1 0 8280 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_185
timestamp 18001
transform 1 0 13432 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_186
timestamp 18001
transform 1 0 18584 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_187
timestamp 18001
transform 1 0 23736 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_188
timestamp 18001
transform 1 0 28888 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_189
timestamp 18001
transform 1 0 5704 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_190
timestamp 18001
transform 1 0 10856 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_191
timestamp 18001
transform 1 0 16008 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_192
timestamp 18001
transform 1 0 21160 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_193
timestamp 18001
transform 1 0 26312 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_194
timestamp 18001
transform 1 0 3128 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_195
timestamp 18001
transform 1 0 8280 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_196
timestamp 18001
transform 1 0 13432 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_197
timestamp 18001
transform 1 0 18584 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_198
timestamp 18001
transform 1 0 23736 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_199
timestamp 18001
transform 1 0 28888 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_200
timestamp 18001
transform 1 0 5704 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_201
timestamp 18001
transform 1 0 10856 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_202
timestamp 18001
transform 1 0 16008 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_203
timestamp 18001
transform 1 0 21160 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_204
timestamp 18001
transform 1 0 26312 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_205
timestamp 18001
transform 1 0 3128 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_206
timestamp 18001
transform 1 0 8280 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_207
timestamp 18001
transform 1 0 13432 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_208
timestamp 18001
transform 1 0 18584 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_209
timestamp 18001
transform 1 0 23736 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_210
timestamp 18001
transform 1 0 28888 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_211
timestamp 18001
transform 1 0 5704 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_212
timestamp 18001
transform 1 0 10856 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_213
timestamp 18001
transform 1 0 16008 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_214
timestamp 18001
transform 1 0 21160 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_215
timestamp 18001
transform 1 0 26312 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_216
timestamp 18001
transform 1 0 3128 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_217
timestamp 18001
transform 1 0 8280 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_218
timestamp 18001
transform 1 0 13432 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_219
timestamp 18001
transform 1 0 18584 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_220
timestamp 18001
transform 1 0 23736 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_221
timestamp 18001
transform 1 0 28888 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_222
timestamp 18001
transform 1 0 5704 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_223
timestamp 18001
transform 1 0 10856 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_224
timestamp 18001
transform 1 0 16008 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_225
timestamp 18001
transform 1 0 21160 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_226
timestamp 18001
transform 1 0 26312 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_227
timestamp 18001
transform 1 0 3128 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_228
timestamp 18001
transform 1 0 8280 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_229
timestamp 18001
transform 1 0 13432 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_230
timestamp 18001
transform 1 0 18584 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_231
timestamp 18001
transform 1 0 23736 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_232
timestamp 18001
transform 1 0 28888 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_233
timestamp 18001
transform 1 0 5704 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_234
timestamp 18001
transform 1 0 10856 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_235
timestamp 18001
transform 1 0 16008 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_236
timestamp 18001
transform 1 0 21160 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_237
timestamp 18001
transform 1 0 26312 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_238
timestamp 18001
transform 1 0 3128 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_239
timestamp 18001
transform 1 0 8280 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_240
timestamp 18001
transform 1 0 13432 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_241
timestamp 18001
transform 1 0 18584 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_242
timestamp 18001
transform 1 0 23736 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_243
timestamp 18001
transform 1 0 28888 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_244
timestamp 18001
transform 1 0 5704 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_245
timestamp 18001
transform 1 0 10856 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_246
timestamp 18001
transform 1 0 16008 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_247
timestamp 18001
transform 1 0 21160 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_248
timestamp 18001
transform 1 0 26312 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_249
timestamp 18001
transform 1 0 3128 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_250
timestamp 18001
transform 1 0 8280 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_251
timestamp 18001
transform 1 0 13432 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_252
timestamp 18001
transform 1 0 18584 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_253
timestamp 18001
transform 1 0 23736 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_254
timestamp 18001
transform 1 0 28888 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_255
timestamp 18001
transform 1 0 3128 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_256
timestamp 18001
transform 1 0 5704 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_257
timestamp 18001
transform 1 0 8280 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_258
timestamp 18001
transform 1 0 10856 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_259
timestamp 18001
transform 1 0 13432 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_260
timestamp 18001
transform 1 0 16008 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_261
timestamp 18001
transform 1 0 18584 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_262
timestamp 18001
transform 1 0 21160 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_263
timestamp 18001
transform 1 0 23736 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_264
timestamp 18001
transform 1 0 26312 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_265
timestamp 18001
transform 1 0 28888 0 -1 19040
box -38 -48 130 592
<< labels >>
flabel metal4 s 4316 496 4636 19088 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 12090 496 12410 19088 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 19864 496 20184 19088 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 27638 496 27958 19088 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 3656 496 3976 19088 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 11430 496 11750 19088 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 19204 496 19524 19088 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 26978 496 27298 19088 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 16118 0 16174 400 0 FreeSans 224 90 0 0 clk
port 2 nsew signal input
flabel metal2 s 18 0 74 400 0 FreeSans 224 90 0 0 ena
port 3 nsew signal input
flabel metal2 s 16762 0 16818 400 0 FreeSans 224 90 0 0 rst_n
port 4 nsew signal input
flabel metal2 s 14186 19600 14242 20000 0 FreeSans 224 90 0 0 ui_in[0]
port 5 nsew signal input
flabel metal2 s 1950 0 2006 400 0 FreeSans 224 90 0 0 ui_in[1]
port 6 nsew signal input
flabel metal2 s 1306 0 1362 400 0 FreeSans 224 90 0 0 ui_in[2]
port 7 nsew signal input
flabel metal2 s 3238 0 3294 400 0 FreeSans 224 90 0 0 ui_in[3]
port 8 nsew signal input
flabel metal2 s 2594 0 2650 400 0 FreeSans 224 90 0 0 ui_in[4]
port 9 nsew signal input
flabel metal2 s 4526 0 4582 400 0 FreeSans 224 90 0 0 ui_in[5]
port 10 nsew signal input
flabel metal2 s 3882 0 3938 400 0 FreeSans 224 90 0 0 ui_in[6]
port 11 nsew signal input
flabel metal2 s 5814 0 5870 400 0 FreeSans 224 90 0 0 ui_in[7]
port 12 nsew signal input
flabel metal2 s 5170 0 5226 400 0 FreeSans 224 90 0 0 uio_in[0]
port 13 nsew signal input
flabel metal2 s 7746 0 7802 400 0 FreeSans 224 90 0 0 uio_in[1]
port 14 nsew signal input
flabel metal2 s 6458 0 6514 400 0 FreeSans 224 90 0 0 uio_in[2]
port 15 nsew signal input
flabel metal2 s 10322 0 10378 400 0 FreeSans 224 90 0 0 uio_in[3]
port 16 nsew signal input
flabel metal2 s 10966 0 11022 400 0 FreeSans 224 90 0 0 uio_in[4]
port 17 nsew signal input
flabel metal2 s 8390 0 8446 400 0 FreeSans 224 90 0 0 uio_in[5]
port 18 nsew signal input
flabel metal2 s 662 0 718 400 0 FreeSans 224 90 0 0 uio_in[6]
port 19 nsew signal input
flabel metal2 s 9678 0 9734 400 0 FreeSans 224 90 0 0 uio_in[7]
port 20 nsew signal input
flabel metal2 s 17406 0 17462 400 0 FreeSans 224 90 0 0 uio_oe[0]
port 21 nsew signal output
flabel metal2 s 18694 0 18750 400 0 FreeSans 224 90 0 0 uio_oe[1]
port 22 nsew signal output
flabel metal2 s 11610 0 11666 400 0 FreeSans 224 90 0 0 uio_oe[2]
port 23 nsew signal output
flabel metal2 s 12254 19600 12310 20000 0 FreeSans 224 90 0 0 uio_oe[3]
port 24 nsew signal output
flabel metal2 s 13542 19600 13598 20000 0 FreeSans 224 90 0 0 uio_oe[4]
port 25 nsew signal output
flabel metal2 s 13542 0 13598 400 0 FreeSans 224 90 0 0 uio_oe[5]
port 26 nsew signal output
flabel metal3 s 0 18368 400 18488 0 FreeSans 480 0 0 0 uio_oe[6]
port 27 nsew signal output
flabel metal2 s 14186 0 14242 400 0 FreeSans 224 90 0 0 uio_oe[7]
port 28 nsew signal output
flabel metal2 s 12254 0 12310 400 0 FreeSans 224 90 0 0 uio_out[0]
port 29 nsew signal output
flabel metal2 s 19982 0 20038 400 0 FreeSans 224 90 0 0 uio_out[1]
port 30 nsew signal output
flabel metal2 s 10322 19600 10378 20000 0 FreeSans 224 90 0 0 uio_out[2]
port 31 nsew signal output
flabel metal2 s 15474 0 15530 400 0 FreeSans 224 90 0 0 uio_out[3]
port 32 nsew signal output
flabel metal3 s 31600 14288 32000 14408 0 FreeSans 480 0 0 0 uio_out[4]
port 33 nsew signal output
flabel metal2 s 7102 0 7158 400 0 FreeSans 224 90 0 0 uio_out[5]
port 34 nsew signal output
flabel metal2 s 9034 0 9090 400 0 FreeSans 224 90 0 0 uio_out[6]
port 35 nsew signal output
flabel metal2 s 16762 19600 16818 20000 0 FreeSans 224 90 0 0 uio_out[7]
port 36 nsew signal output
flabel metal2 s 16118 19600 16174 20000 0 FreeSans 224 90 0 0 uo_out[0]
port 37 nsew signal output
flabel metal2 s 17406 19600 17462 20000 0 FreeSans 224 90 0 0 uo_out[1]
port 38 nsew signal output
flabel metal2 s 14830 19600 14886 20000 0 FreeSans 224 90 0 0 uo_out[2]
port 39 nsew signal output
flabel metal2 s 22558 19600 22614 20000 0 FreeSans 224 90 0 0 uo_out[3]
port 40 nsew signal output
flabel metal2 s 12898 19600 12954 20000 0 FreeSans 224 90 0 0 uo_out[4]
port 41 nsew signal output
flabel metal2 s 18050 0 18106 400 0 FreeSans 224 90 0 0 uo_out[5]
port 42 nsew signal output
flabel metal2 s 14830 0 14886 400 0 FreeSans 224 90 0 0 uo_out[6]
port 43 nsew signal output
flabel metal2 s 12898 0 12954 400 0 FreeSans 224 90 0 0 uo_out[7]
port 44 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 32000 20000
<< end >>
