magic
tech sky130A
magscale 1 2
timestamp 1768779796
<< viali >>
rect 11805 28713 11839 28747
rect 12449 28713 12483 28747
rect 13093 28713 13127 28747
rect 13737 28713 13771 28747
rect 14381 28713 14415 28747
rect 15025 28713 15059 28747
rect 15669 28713 15703 28747
rect 16313 28713 16347 28747
rect 16957 28713 16991 28747
rect 17601 28713 17635 28747
rect 18245 28713 18279 28747
rect 18889 28713 18923 28747
rect 19625 28713 19659 28747
rect 20269 28713 20303 28747
rect 20913 28713 20947 28747
rect 21557 28713 21591 28747
rect 22109 28713 22143 28747
rect 22845 28713 22879 28747
rect 23489 28713 23523 28747
rect 24133 28713 24167 28747
rect 24777 28713 24811 28747
rect 25421 28713 25455 28747
rect 26065 28713 26099 28747
rect 26709 28713 26743 28747
rect 27353 28713 27387 28747
rect 27721 28713 27755 28747
rect 11989 28509 12023 28543
rect 12633 28509 12667 28543
rect 13277 28509 13311 28543
rect 13921 28509 13955 28543
rect 14565 28509 14599 28543
rect 15209 28509 15243 28543
rect 15853 28509 15887 28543
rect 16497 28509 16531 28543
rect 17141 28509 17175 28543
rect 17785 28509 17819 28543
rect 18429 28509 18463 28543
rect 19073 28509 19107 28543
rect 19441 28509 19475 28543
rect 20085 28509 20119 28543
rect 20729 28509 20763 28543
rect 21373 28509 21407 28543
rect 22293 28509 22327 28543
rect 22661 28509 22695 28543
rect 23305 28509 23339 28543
rect 23949 28509 23983 28543
rect 24593 28509 24627 28543
rect 25237 28509 25271 28543
rect 25881 28509 25915 28543
rect 26525 28509 26559 28543
rect 27169 28509 27203 28543
rect 27537 28509 27571 28543
rect 18981 28169 19015 28203
rect 20177 28169 20211 28203
rect 20453 28169 20487 28203
rect 24961 28169 24995 28203
rect 27721 28169 27755 28203
rect 19625 28101 19659 28135
rect 11099 28033 11133 28067
rect 11253 28033 11287 28067
rect 18705 28033 18739 28067
rect 19165 28033 19199 28067
rect 19257 28033 19291 28067
rect 19349 28033 19383 28067
rect 19809 28033 19843 28067
rect 20091 28033 20125 28067
rect 20269 28033 20303 28067
rect 20361 28033 20395 28067
rect 20545 28033 20579 28067
rect 21649 28033 21683 28067
rect 22017 28033 22051 28067
rect 22201 28033 22235 28067
rect 24869 28033 24903 28067
rect 25053 28033 25087 28067
rect 27169 28033 27203 28067
rect 27537 28033 27571 28067
rect 10333 27965 10367 27999
rect 19993 27965 20027 27999
rect 10701 27897 10735 27931
rect 10793 27897 10827 27931
rect 19533 27897 19567 27931
rect 27353 27897 27387 27931
rect 11069 27829 11103 27863
rect 18613 27829 18647 27863
rect 21557 27829 21591 27863
rect 22201 27829 22235 27863
rect 6837 27625 6871 27659
rect 10333 27625 10367 27659
rect 18153 27625 18187 27659
rect 18797 27625 18831 27659
rect 19901 27625 19935 27659
rect 20085 27625 20119 27659
rect 20821 27625 20855 27659
rect 21373 27625 21407 27659
rect 22385 27625 22419 27659
rect 23765 27625 23799 27659
rect 24225 27625 24259 27659
rect 24869 27625 24903 27659
rect 25145 27625 25179 27659
rect 25697 27625 25731 27659
rect 26157 27625 26191 27659
rect 26801 27625 26835 27659
rect 27261 27625 27295 27659
rect 10701 27557 10735 27591
rect 16957 27557 16991 27591
rect 17233 27557 17267 27591
rect 18613 27557 18647 27591
rect 21097 27557 21131 27591
rect 21465 27557 21499 27591
rect 22201 27557 22235 27591
rect 5089 27489 5123 27523
rect 5276 27489 5310 27523
rect 6653 27489 6687 27523
rect 7021 27489 7055 27523
rect 17509 27489 17543 27523
rect 21741 27489 21775 27523
rect 22753 27489 22787 27523
rect 24501 27489 24535 27523
rect 25311 27489 25345 27523
rect 26341 27489 26375 27523
rect 4997 27421 5031 27455
rect 5365 27421 5399 27455
rect 5549 27421 5583 27455
rect 5825 27421 5859 27455
rect 6009 27421 6043 27455
rect 6101 27421 6135 27455
rect 6193 27421 6227 27455
rect 6285 27421 6319 27455
rect 6561 27421 6595 27455
rect 7205 27399 7239 27433
rect 7481 27421 7515 27455
rect 7665 27421 7699 27455
rect 9505 27421 9539 27455
rect 9965 27421 9999 27455
rect 10333 27421 10367 27455
rect 10609 27421 10643 27455
rect 10793 27421 10827 27455
rect 11161 27421 11195 27455
rect 11437 27421 11471 27455
rect 11743 27421 11777 27455
rect 11897 27421 11931 27455
rect 16957 27421 16991 27455
rect 17141 27421 17175 27455
rect 17233 27421 17267 27455
rect 17417 27421 17451 27455
rect 17784 27421 17818 27455
rect 17877 27421 17911 27455
rect 18521 27421 18555 27455
rect 19441 27421 19475 27455
rect 19533 27421 19567 27455
rect 20453 27421 20487 27455
rect 20545 27421 20579 27455
rect 20913 27421 20947 27455
rect 21189 27421 21223 27455
rect 21373 27421 21407 27455
rect 23029 27421 23063 27455
rect 23121 27421 23155 27455
rect 23397 27421 23431 27455
rect 24041 27421 24075 27455
rect 24225 27421 24259 27455
rect 24593 27421 24627 27455
rect 24961 27421 24995 27455
rect 25421 27421 25455 27455
rect 25789 27421 25823 27455
rect 26065 27421 26099 27455
rect 26525 27421 26559 27455
rect 26801 27421 26835 27455
rect 26985 27421 27019 27455
rect 27077 27421 27111 27455
rect 27261 27421 27295 27455
rect 9689 27353 9723 27387
rect 9873 27353 9907 27387
rect 18981 27353 19015 27387
rect 19809 27353 19843 27387
rect 21649 27353 21683 27387
rect 22201 27353 22235 27387
rect 22544 27353 22578 27387
rect 22661 27353 22695 27387
rect 23489 27353 23523 27387
rect 23606 27353 23640 27387
rect 5273 27285 5307 27319
rect 5457 27285 5491 27319
rect 5825 27285 5859 27319
rect 10517 27285 10551 27319
rect 11529 27285 11563 27319
rect 17969 27285 18003 27319
rect 18153 27285 18187 27319
rect 18771 27285 18805 27319
rect 19257 27285 19291 27319
rect 19625 27285 19659 27319
rect 20085 27285 20119 27319
rect 25973 27285 26007 27319
rect 26709 27285 26743 27319
rect 5089 27081 5123 27115
rect 5983 27081 6017 27115
rect 11253 27081 11287 27115
rect 12541 27081 12575 27115
rect 17417 27081 17451 27115
rect 18153 27081 18187 27115
rect 18705 27081 18739 27115
rect 19625 27081 19659 27115
rect 21005 27081 21039 27115
rect 22201 27081 22235 27115
rect 22385 27081 22419 27115
rect 23213 27081 23247 27115
rect 24777 27081 24811 27115
rect 24961 27081 24995 27115
rect 25973 27081 26007 27115
rect 2789 27013 2823 27047
rect 2989 27013 3023 27047
rect 6193 27013 6227 27047
rect 11681 27013 11715 27047
rect 11897 27013 11931 27047
rect 11989 27013 12023 27047
rect 12173 27013 12207 27047
rect 18305 27013 18339 27047
rect 18521 27013 18555 27047
rect 21097 27013 21131 27047
rect 22017 27013 22051 27047
rect 25421 27013 25455 27047
rect 2237 26945 2271 26979
rect 3525 26945 3559 26979
rect 3709 26945 3743 26979
rect 3985 26945 4019 26979
rect 4721 26945 4755 26979
rect 5365 26945 5399 26979
rect 5549 26945 5583 26979
rect 6561 26945 6595 26979
rect 7021 26945 7055 26979
rect 7113 26945 7147 26979
rect 7389 26945 7423 26979
rect 9137 26945 9171 26979
rect 10701 26945 10735 26979
rect 10793 26945 10827 26979
rect 10977 26945 11011 26979
rect 11161 26945 11195 26979
rect 12357 26945 12391 26979
rect 12449 26945 12483 26979
rect 12725 26945 12759 26979
rect 17325 26945 17359 26979
rect 17509 26945 17543 26979
rect 17877 26945 17911 26979
rect 18061 26945 18095 26979
rect 18613 26945 18647 26979
rect 18797 26945 18831 26979
rect 19073 26945 19107 26979
rect 19533 26945 19567 26979
rect 19809 26945 19843 26979
rect 20269 26945 20303 26979
rect 20361 26945 20395 26979
rect 20545 26945 20579 26979
rect 20821 26945 20855 26979
rect 21311 26945 21345 26979
rect 21465 26945 21499 26979
rect 22109 26945 22143 26979
rect 22661 26945 22695 26979
rect 22937 26945 22971 26979
rect 23029 26945 23063 26979
rect 24133 26945 24167 26979
rect 24593 26945 24627 26979
rect 24869 26945 24903 26979
rect 25053 26945 25087 26979
rect 25329 26945 25363 26979
rect 25513 26945 25547 26979
rect 25881 26945 25915 26979
rect 26065 26945 26099 26979
rect 26157 26945 26191 26979
rect 26341 26945 26375 26979
rect 2145 26877 2179 26911
rect 2605 26877 2639 26911
rect 3249 26877 3283 26911
rect 3893 26877 3927 26911
rect 4813 26877 4847 26911
rect 5273 26877 5307 26911
rect 5457 26877 5491 26911
rect 5733 26877 5767 26911
rect 7205 26877 7239 26911
rect 9229 26877 9263 26911
rect 9781 26877 9815 26911
rect 9873 26877 9907 26911
rect 10241 26877 10275 26911
rect 10885 26877 10919 26911
rect 19165 26877 19199 26911
rect 19993 26877 20027 26911
rect 20729 26877 20763 26911
rect 22569 26877 22603 26911
rect 24501 26877 24535 26911
rect 3525 26809 3559 26843
rect 5825 26809 5859 26843
rect 6699 26809 6733 26843
rect 17877 26809 17911 26843
rect 18889 26809 18923 26843
rect 20637 26809 20671 26843
rect 21833 26809 21867 26843
rect 26157 26809 26191 26843
rect 2973 26741 3007 26775
rect 3157 26741 3191 26775
rect 4261 26741 4295 26775
rect 6009 26741 6043 26775
rect 6837 26741 6871 26775
rect 6929 26741 6963 26775
rect 7113 26741 7147 26775
rect 7573 26741 7607 26775
rect 8861 26741 8895 26775
rect 9597 26741 9631 26775
rect 10517 26741 10551 26775
rect 11529 26741 11563 26775
rect 11713 26741 11747 26775
rect 12725 26741 12759 26775
rect 18337 26741 18371 26775
rect 19073 26741 19107 26775
rect 20177 26741 20211 26775
rect 24225 26741 24259 26775
rect 3985 26537 4019 26571
rect 5457 26537 5491 26571
rect 7021 26537 7055 26571
rect 10701 26537 10735 26571
rect 11069 26537 11103 26571
rect 19441 26537 19475 26571
rect 19625 26537 19659 26571
rect 22845 26537 22879 26571
rect 25053 26537 25087 26571
rect 26065 26537 26099 26571
rect 26709 26537 26743 26571
rect 3157 26469 3191 26503
rect 27721 26469 27755 26503
rect 6285 26401 6319 26435
rect 6745 26401 6779 26435
rect 20085 26401 20119 26435
rect 25145 26401 25179 26435
rect 25630 26401 25664 26435
rect 1777 26333 1811 26367
rect 2881 26333 2915 26367
rect 3157 26333 3191 26367
rect 3801 26333 3835 26367
rect 3985 26333 4019 26367
rect 4997 26333 5031 26367
rect 5273 26333 5307 26367
rect 5365 26333 5399 26367
rect 5549 26333 5583 26367
rect 5641 26333 5675 26367
rect 5825 26333 5859 26367
rect 6193 26333 6227 26367
rect 6653 26333 6687 26367
rect 6837 26333 6871 26367
rect 7113 26333 7147 26367
rect 7481 26333 7515 26367
rect 7665 26333 7699 26367
rect 8493 26333 8527 26367
rect 8585 26333 8619 26367
rect 8769 26333 8803 26367
rect 8953 26333 8987 26367
rect 9045 26333 9079 26367
rect 9229 26333 9263 26367
rect 9781 26333 9815 26367
rect 10057 26333 10091 26367
rect 10333 26333 10367 26367
rect 10517 26333 10551 26367
rect 10609 26333 10643 26367
rect 10885 26333 10919 26367
rect 11161 26333 11195 26367
rect 12265 26333 12299 26367
rect 12541 26333 12575 26367
rect 12817 26333 12851 26367
rect 13093 26333 13127 26367
rect 13185 26333 13219 26367
rect 13277 26333 13311 26367
rect 13461 26333 13495 26367
rect 19993 26333 20027 26367
rect 20269 26333 20303 26367
rect 20453 26333 20487 26367
rect 20913 26333 20947 26367
rect 21005 26333 21039 26367
rect 23121 26333 23155 26367
rect 24869 26333 24903 26367
rect 25513 26333 25547 26367
rect 26525 26333 26559 26367
rect 26709 26333 26743 26367
rect 27537 26333 27571 26367
rect 2513 26265 2547 26299
rect 5089 26265 5123 26299
rect 5733 26265 5767 26299
rect 9965 26265 9999 26299
rect 12081 26265 12115 26299
rect 22937 26265 22971 26299
rect 26157 26265 26191 26299
rect 26341 26265 26375 26299
rect 2973 26197 3007 26231
rect 5174 26197 5208 26231
rect 6561 26197 6595 26231
rect 7665 26197 7699 26231
rect 8677 26197 8711 26231
rect 9413 26197 9447 26231
rect 10057 26197 10091 26231
rect 10149 26197 10183 26231
rect 12449 26197 12483 26231
rect 12633 26197 12667 26231
rect 13001 26197 13035 26231
rect 13185 26197 13219 26231
rect 19625 26197 19659 26231
rect 25421 26197 25455 26231
rect 25789 26197 25823 26231
rect 2789 25993 2823 26027
rect 8125 25993 8159 26027
rect 12725 25993 12759 26027
rect 26449 25993 26483 26027
rect 26617 25993 26651 26027
rect 7757 25925 7791 25959
rect 26249 25925 26283 25959
rect 3065 25857 3099 25891
rect 7941 25857 7975 25891
rect 10425 25857 10459 25891
rect 10609 25857 10643 25891
rect 12541 25857 12575 25891
rect 12725 25857 12759 25891
rect 26985 25857 27019 25891
rect 10517 25653 10551 25687
rect 26433 25653 26467 25687
rect 27077 25653 27111 25687
rect 20453 25449 20487 25483
rect 20637 25449 20671 25483
rect 21005 25449 21039 25483
rect 23397 25449 23431 25483
rect 27169 25449 27203 25483
rect 7205 25381 7239 25415
rect 22937 25381 22971 25415
rect 26341 25381 26375 25415
rect 2513 25313 2547 25347
rect 6561 25313 6595 25347
rect 6929 25313 6963 25347
rect 7665 25313 7699 25347
rect 15117 25313 15151 25347
rect 26157 25313 26191 25347
rect 2789 25245 2823 25279
rect 6469 25245 6503 25279
rect 7573 25245 7607 25279
rect 7757 25245 7791 25279
rect 8033 25245 8067 25279
rect 8217 25245 8251 25279
rect 9321 25245 9355 25279
rect 9505 25245 9539 25279
rect 10057 25245 10091 25279
rect 10211 25245 10245 25279
rect 12357 25245 12391 25279
rect 12449 25245 12483 25279
rect 12633 25245 12667 25279
rect 12725 25245 12759 25279
rect 15485 25245 15519 25279
rect 15577 25245 15611 25279
rect 15945 25245 15979 25279
rect 16037 25245 16071 25279
rect 16129 25245 16163 25279
rect 21097 25245 21131 25279
rect 22477 25245 22511 25279
rect 22661 25245 22695 25279
rect 22845 25245 22879 25279
rect 23213 25245 23247 25279
rect 25789 25245 25823 25279
rect 25881 25245 25915 25279
rect 26249 25245 26283 25279
rect 26525 25245 26559 25279
rect 27537 25245 27571 25279
rect 15761 25177 15795 25211
rect 20821 25177 20855 25211
rect 22937 25177 22971 25211
rect 23121 25177 23155 25211
rect 23489 25177 23523 25211
rect 25605 25177 25639 25211
rect 25973 25177 26007 25211
rect 26709 25177 26743 25211
rect 26801 25177 26835 25211
rect 26985 25177 27019 25211
rect 3433 25109 3467 25143
rect 6837 25109 6871 25143
rect 7389 25109 7423 25143
rect 8217 25109 8251 25143
rect 9505 25109 9539 25143
rect 10425 25109 10459 25143
rect 12909 25109 12943 25143
rect 16313 25109 16347 25143
rect 20621 25109 20655 25143
rect 27721 25109 27755 25143
rect 12081 24905 12115 24939
rect 17433 24905 17467 24939
rect 10057 24837 10091 24871
rect 12909 24837 12943 24871
rect 17233 24837 17267 24871
rect 26157 24837 26191 24871
rect 4261 24769 4295 24803
rect 7941 24769 7975 24803
rect 8125 24769 8159 24803
rect 8401 24769 8435 24803
rect 8769 24769 8803 24803
rect 9873 24769 9907 24803
rect 10333 24769 10367 24803
rect 10517 24769 10551 24803
rect 10609 24769 10643 24803
rect 10701 24769 10735 24803
rect 11805 24769 11839 24803
rect 12173 24769 12207 24803
rect 12265 24769 12299 24803
rect 12725 24769 12759 24803
rect 13001 24769 13035 24803
rect 13185 24769 13219 24803
rect 15025 24769 15059 24803
rect 15117 24769 15151 24803
rect 15301 24769 15335 24803
rect 15577 24769 15611 24803
rect 15761 24769 15795 24803
rect 15853 24769 15887 24803
rect 16313 24769 16347 24803
rect 16497 24769 16531 24803
rect 16681 24769 16715 24803
rect 16773 24769 16807 24803
rect 16957 24769 16991 24803
rect 21925 24769 21959 24803
rect 22293 24769 22327 24803
rect 25237 24769 25271 24803
rect 25513 24769 25547 24803
rect 26617 24769 26651 24803
rect 26985 24769 27019 24803
rect 27077 24769 27111 24803
rect 27169 24769 27203 24803
rect 27537 24769 27571 24803
rect 4169 24701 4203 24735
rect 4353 24701 4387 24735
rect 4445 24701 4479 24735
rect 8861 24701 8895 24735
rect 8953 24701 8987 24735
rect 10977 24701 11011 24735
rect 11621 24701 11655 24735
rect 12541 24701 12575 24735
rect 17141 24701 17175 24735
rect 22201 24701 22235 24735
rect 22569 24701 22603 24735
rect 24041 24701 24075 24735
rect 25421 24701 25455 24735
rect 26065 24701 26099 24735
rect 26525 24701 26559 24735
rect 12357 24633 12391 24667
rect 22017 24633 22051 24667
rect 25513 24633 25547 24667
rect 25789 24633 25823 24667
rect 26801 24633 26835 24667
rect 4629 24565 4663 24599
rect 8585 24565 8619 24599
rect 9137 24565 9171 24599
rect 10241 24565 10275 24599
rect 12449 24565 12483 24599
rect 13185 24565 13219 24599
rect 15485 24565 15519 24599
rect 15853 24565 15887 24599
rect 16405 24565 16439 24599
rect 17417 24565 17451 24599
rect 17601 24565 17635 24599
rect 22109 24565 22143 24599
rect 25605 24565 25639 24599
rect 26249 24565 26283 24599
rect 27721 24565 27755 24599
rect 3617 24361 3651 24395
rect 5365 24361 5399 24395
rect 7573 24361 7607 24395
rect 11989 24361 12023 24395
rect 12173 24361 12207 24395
rect 21005 24361 21039 24395
rect 21741 24361 21775 24395
rect 23857 24361 23891 24395
rect 24041 24361 24075 24395
rect 26341 24361 26375 24395
rect 26433 24361 26467 24395
rect 27261 24361 27295 24395
rect 9321 24293 9355 24327
rect 10149 24293 10183 24327
rect 10517 24293 10551 24327
rect 24409 24293 24443 24327
rect 27445 24293 27479 24327
rect 7205 24225 7239 24259
rect 9965 24225 9999 24259
rect 13737 24225 13771 24259
rect 15301 24225 15335 24259
rect 18153 24225 18187 24259
rect 19257 24225 19291 24259
rect 21833 24225 21867 24259
rect 21925 24225 21959 24259
rect 24961 24225 24995 24259
rect 25145 24225 25179 24259
rect 25605 24225 25639 24259
rect 26985 24225 27019 24259
rect 1409 24157 1443 24191
rect 1777 24157 1811 24191
rect 2881 24157 2915 24191
rect 3065 24157 3099 24191
rect 3433 24157 3467 24191
rect 3617 24157 3651 24191
rect 3893 24157 3927 24191
rect 4997 24157 5031 24191
rect 5181 24157 5215 24191
rect 5273 24157 5307 24191
rect 7389 24157 7423 24191
rect 9137 24157 9171 24191
rect 9403 24157 9437 24191
rect 9505 24157 9539 24191
rect 9689 24157 9723 24191
rect 9781 24157 9815 24191
rect 10057 24157 10091 24191
rect 10333 24157 10367 24191
rect 10425 24157 10459 24191
rect 12633 24157 12667 24191
rect 12909 24157 12943 24191
rect 13001 24157 13035 24191
rect 13369 24157 13403 24191
rect 14105 24157 14139 24191
rect 14289 24157 14323 24191
rect 17325 24157 17359 24191
rect 17555 24157 17589 24191
rect 17693 24157 17727 24191
rect 17785 24157 17819 24191
rect 18245 24157 18279 24191
rect 21557 24157 21591 24191
rect 24685 24157 24719 24191
rect 25237 24157 25271 24191
rect 25697 24157 25731 24191
rect 25845 24157 25879 24191
rect 26203 24157 26237 24191
rect 26617 24157 26651 24191
rect 27537 24157 27571 24191
rect 2513 24089 2547 24123
rect 2973 24089 3007 24123
rect 4629 24089 4663 24123
rect 8953 24089 8987 24123
rect 11805 24089 11839 24123
rect 12021 24089 12055 24123
rect 15577 24089 15611 24123
rect 17417 24089 17451 24123
rect 19533 24089 19567 24123
rect 22201 24089 22235 24123
rect 24025 24089 24059 24123
rect 24225 24089 24259 24123
rect 24409 24089 24443 24123
rect 25513 24089 25547 24123
rect 25973 24089 26007 24123
rect 26065 24089 26099 24123
rect 27077 24089 27111 24123
rect 27277 24089 27311 24123
rect 1593 24021 1627 24055
rect 5181 24021 5215 24055
rect 14473 24021 14507 24055
rect 17049 24021 17083 24055
rect 17141 24021 17175 24055
rect 17877 24021 17911 24055
rect 21373 24021 21407 24055
rect 23673 24021 23707 24055
rect 24593 24021 24627 24055
rect 25421 24021 25455 24055
rect 26801 24021 26835 24055
rect 27721 24021 27755 24055
rect 8953 23817 8987 23851
rect 9873 23817 9907 23851
rect 16865 23817 16899 23851
rect 17509 23817 17543 23851
rect 17601 23817 17635 23851
rect 17985 23817 18019 23851
rect 18981 23817 19015 23851
rect 23765 23817 23799 23851
rect 25421 23817 25455 23851
rect 3157 23749 3191 23783
rect 9505 23749 9539 23783
rect 16773 23749 16807 23783
rect 17785 23749 17819 23783
rect 22109 23749 22143 23783
rect 25513 23749 25547 23783
rect 1501 23681 1535 23715
rect 2421 23681 2455 23715
rect 2513 23681 2547 23715
rect 3525 23681 3559 23715
rect 4353 23681 4387 23715
rect 5273 23681 5307 23715
rect 8861 23681 8895 23715
rect 9045 23681 9079 23715
rect 9689 23681 9723 23715
rect 12081 23681 12115 23715
rect 12265 23681 12299 23715
rect 12449 23681 12483 23715
rect 12633 23681 12667 23715
rect 13185 23681 13219 23715
rect 15761 23681 15795 23715
rect 15945 23681 15979 23715
rect 16497 23681 16531 23715
rect 16681 23681 16715 23715
rect 17141 23681 17175 23715
rect 17325 23681 17359 23715
rect 17693 23681 17727 23715
rect 18613 23681 18647 23715
rect 18889 23681 18923 23715
rect 19441 23681 19475 23715
rect 19625 23681 19659 23715
rect 19717 23681 19751 23715
rect 21833 23681 21867 23715
rect 23673 23681 23707 23715
rect 23857 23681 23891 23715
rect 24961 23681 24995 23715
rect 25697 23681 25731 23715
rect 27537 23681 27571 23715
rect 3065 23613 3099 23647
rect 4445 23613 4479 23647
rect 4905 23613 4939 23647
rect 5181 23613 5215 23647
rect 12357 23613 12391 23647
rect 12909 23613 12943 23647
rect 19257 23613 19291 23647
rect 25053 23613 25087 23647
rect 17141 23545 17175 23579
rect 18705 23545 18739 23579
rect 23581 23545 23615 23579
rect 1777 23477 1811 23511
rect 5641 23477 5675 23511
rect 12173 23477 12207 23511
rect 12817 23477 12851 23511
rect 13001 23477 13035 23511
rect 13369 23477 13403 23511
rect 15853 23477 15887 23511
rect 16405 23477 16439 23511
rect 17049 23477 17083 23511
rect 17417 23477 17451 23511
rect 17969 23477 18003 23511
rect 18153 23477 18187 23511
rect 24777 23477 24811 23511
rect 27721 23477 27755 23511
rect 4353 23273 4387 23307
rect 10425 23273 10459 23307
rect 13001 23273 13035 23307
rect 19073 23273 19107 23307
rect 19625 23273 19659 23307
rect 22477 23273 22511 23307
rect 22845 23273 22879 23307
rect 26801 23273 26835 23307
rect 4905 23205 4939 23239
rect 8217 23205 8251 23239
rect 10977 23205 11011 23239
rect 19993 23205 20027 23239
rect 20361 23205 20395 23239
rect 26709 23205 26743 23239
rect 5181 23137 5215 23171
rect 5549 23137 5583 23171
rect 7389 23137 7423 23171
rect 9229 23137 9263 23171
rect 12817 23137 12851 23171
rect 22937 23137 22971 23171
rect 24409 23137 24443 23171
rect 4261 23069 4295 23103
rect 4445 23069 4479 23103
rect 4905 23069 4939 23103
rect 5089 23069 5123 23103
rect 5641 23069 5675 23103
rect 5825 23069 5859 23103
rect 6193 23069 6227 23103
rect 7481 23069 7515 23103
rect 7941 23069 7975 23103
rect 9137 23069 9171 23103
rect 9413 23069 9447 23103
rect 9781 23069 9815 23103
rect 9873 23069 9907 23103
rect 9965 23069 9999 23103
rect 10149 23069 10183 23103
rect 10241 23069 10275 23103
rect 10517 23069 10551 23103
rect 10609 23069 10643 23103
rect 10793 23069 10827 23103
rect 12357 23069 12391 23103
rect 12449 23069 12483 23103
rect 12633 23069 12667 23103
rect 12909 23069 12943 23103
rect 13277 23069 13311 23103
rect 18521 23069 18555 23103
rect 18705 23069 18739 23103
rect 18981 23069 19015 23103
rect 19073 23069 19107 23103
rect 20085 23069 20119 23103
rect 20361 23069 20395 23103
rect 20453 23069 20487 23103
rect 20637 23069 20671 23103
rect 22661 23069 22695 23103
rect 23213 23069 23247 23103
rect 24041 23069 24075 23103
rect 24225 23069 24259 23103
rect 26617 23069 26651 23103
rect 7205 23001 7239 23035
rect 8217 23001 8251 23035
rect 9597 23001 9631 23035
rect 18797 23001 18831 23035
rect 19625 23001 19659 23035
rect 23029 23001 23063 23035
rect 24133 23001 24167 23035
rect 24685 23001 24719 23035
rect 26893 23001 26927 23035
rect 7849 22933 7883 22967
rect 8033 22933 8067 22967
rect 13461 22933 13495 22967
rect 18705 22933 18739 22967
rect 19441 22933 19475 22967
rect 20177 22933 20211 22967
rect 20545 22933 20579 22967
rect 26157 22933 26191 22967
rect 7957 22729 7991 22763
rect 8125 22729 8159 22763
rect 10333 22729 10367 22763
rect 13645 22729 13679 22763
rect 14305 22729 14339 22763
rect 17141 22729 17175 22763
rect 20821 22729 20855 22763
rect 26433 22729 26467 22763
rect 27185 22729 27219 22763
rect 1501 22661 1535 22695
rect 6561 22661 6595 22695
rect 7757 22661 7791 22695
rect 8677 22661 8711 22695
rect 8861 22661 8895 22695
rect 9597 22661 9631 22695
rect 9965 22661 9999 22695
rect 14105 22661 14139 22695
rect 16773 22661 16807 22695
rect 16989 22661 17023 22695
rect 21373 22661 21407 22695
rect 26985 22661 27019 22695
rect 2237 22593 2271 22627
rect 2421 22593 2455 22627
rect 3709 22593 3743 22627
rect 3893 22593 3927 22627
rect 5549 22593 5583 22627
rect 6469 22593 6503 22627
rect 6653 22593 6687 22627
rect 9505 22593 9539 22627
rect 9781 22593 9815 22627
rect 10057 22593 10091 22627
rect 10241 22593 10275 22627
rect 10333 22593 10367 22627
rect 12817 22593 12851 22627
rect 13277 22593 13311 22627
rect 17233 22593 17267 22627
rect 17417 22593 17451 22627
rect 17509 22593 17543 22627
rect 19349 22593 19383 22627
rect 21005 22593 21039 22627
rect 21281 22593 21315 22627
rect 21465 22593 21499 22627
rect 25697 22593 25731 22627
rect 25881 22593 25915 22627
rect 26065 22593 26099 22627
rect 26525 22593 26559 22627
rect 27537 22593 27571 22627
rect 2329 22525 2363 22559
rect 2789 22525 2823 22559
rect 3617 22525 3651 22559
rect 5641 22525 5675 22559
rect 9045 22525 9079 22559
rect 13185 22525 13219 22559
rect 19441 22525 19475 22559
rect 21189 22525 21223 22559
rect 1685 22457 1719 22491
rect 27353 22457 27387 22491
rect 27721 22457 27755 22491
rect 3893 22389 3927 22423
rect 5917 22389 5951 22423
rect 7941 22389 7975 22423
rect 12909 22389 12943 22423
rect 14289 22389 14323 22423
rect 14473 22389 14507 22423
rect 16957 22389 16991 22423
rect 17233 22389 17267 22423
rect 19625 22389 19659 22423
rect 25513 22389 25547 22423
rect 25973 22389 26007 22423
rect 27169 22389 27203 22423
rect 3065 22185 3099 22219
rect 4537 22185 4571 22219
rect 7389 22185 7423 22219
rect 25789 22185 25823 22219
rect 16313 22117 16347 22151
rect 2237 22049 2271 22083
rect 3893 22049 3927 22083
rect 3985 22049 4019 22083
rect 9321 22049 9355 22083
rect 9689 22049 9723 22083
rect 10609 22049 10643 22083
rect 16865 22049 16899 22083
rect 1409 21981 1443 22015
rect 2145 21981 2179 22015
rect 3249 21981 3283 22015
rect 4077 21981 4111 22015
rect 4169 21981 4203 22015
rect 4445 21981 4479 22015
rect 7297 21981 7331 22015
rect 7481 21981 7515 22015
rect 9229 21981 9263 22015
rect 9413 21981 9447 22015
rect 9781 21981 9815 22015
rect 13369 21981 13403 22015
rect 14657 21981 14691 22015
rect 14933 21981 14967 22015
rect 15301 21981 15335 22015
rect 15485 21981 15519 22015
rect 17141 21981 17175 22015
rect 17325 21981 17359 22015
rect 25237 21981 25271 22015
rect 25329 21981 25363 22015
rect 16313 21913 16347 21947
rect 25513 21913 25547 21947
rect 25973 21913 26007 21947
rect 26157 21913 26191 21947
rect 1593 21845 1627 21879
rect 2881 21845 2915 21879
rect 4353 21845 4387 21879
rect 13461 21845 13495 21879
rect 15209 21845 15243 21879
rect 16773 21845 16807 21879
rect 17049 21845 17083 21879
rect 17509 21845 17543 21879
rect 25237 21845 25271 21879
rect 25605 21845 25639 21879
rect 25773 21845 25807 21879
rect 26249 21845 26283 21879
rect 4445 21641 4479 21675
rect 14473 21641 14507 21675
rect 25263 21641 25297 21675
rect 26065 21641 26099 21675
rect 1961 21573 1995 21607
rect 12725 21573 12759 21607
rect 13369 21573 13403 21607
rect 20453 21573 20487 21607
rect 24685 21573 24719 21607
rect 25053 21573 25087 21607
rect 25605 21573 25639 21607
rect 3801 21505 3835 21539
rect 3985 21505 4019 21539
rect 4629 21505 4663 21539
rect 7389 21505 7423 21539
rect 12633 21505 12667 21539
rect 12817 21505 12851 21539
rect 13093 21505 13127 21539
rect 13185 21505 13219 21539
rect 13553 21505 13587 21539
rect 13645 21503 13679 21537
rect 13921 21505 13955 21539
rect 14289 21505 14323 21539
rect 14933 21505 14967 21539
rect 15117 21505 15151 21539
rect 16129 21505 16163 21539
rect 16313 21505 16347 21539
rect 17141 21505 17175 21539
rect 17601 21505 17635 21539
rect 18061 21505 18095 21539
rect 18429 21505 18463 21539
rect 18981 21505 19015 21539
rect 19625 21505 19659 21539
rect 20545 21505 20579 21539
rect 23121 21505 23155 21539
rect 24869 21505 24903 21539
rect 24961 21505 24995 21539
rect 25513 21505 25547 21539
rect 25789 21505 25823 21539
rect 27169 21505 27203 21539
rect 2513 21437 2547 21471
rect 5641 21437 5675 21471
rect 7297 21437 7331 21471
rect 8125 21437 8159 21471
rect 15301 21437 15335 21471
rect 16221 21437 16255 21471
rect 16497 21437 16531 21471
rect 26525 21437 26559 21471
rect 13829 21369 13863 21403
rect 17233 21369 17267 21403
rect 24685 21369 24719 21403
rect 25421 21369 25455 21403
rect 26157 21369 26191 21403
rect 26985 21369 27019 21403
rect 12909 21301 12943 21335
rect 13369 21301 13403 21335
rect 14289 21301 14323 21335
rect 19809 21301 19843 21335
rect 22845 21301 22879 21335
rect 25237 21301 25271 21335
rect 25973 21301 26007 21335
rect 3893 21097 3927 21131
rect 12357 21097 12391 21131
rect 12817 21097 12851 21131
rect 16497 21097 16531 21131
rect 17141 21097 17175 21131
rect 23581 21097 23615 21131
rect 25053 21097 25087 21131
rect 27077 21097 27111 21131
rect 19533 21029 19567 21063
rect 19625 21029 19659 21063
rect 23121 21029 23155 21063
rect 6377 20961 6411 20995
rect 6837 20961 6871 20995
rect 13001 20961 13035 20995
rect 15209 20961 15243 20995
rect 16681 20961 16715 20995
rect 17325 20961 17359 20995
rect 17417 20961 17451 20995
rect 17693 20961 17727 20995
rect 17785 20961 17819 20995
rect 21557 20961 21591 20995
rect 21741 20961 21775 20995
rect 22569 20961 22603 20995
rect 25605 20961 25639 20995
rect 1961 20893 1995 20927
rect 3801 20893 3835 20927
rect 3985 20893 4019 20927
rect 4813 20893 4847 20927
rect 4997 20893 5031 20927
rect 5641 20893 5675 20927
rect 5733 20893 5767 20927
rect 5917 20893 5951 20927
rect 6469 20893 6503 20927
rect 6929 20893 6963 20927
rect 7113 20893 7147 20927
rect 10609 20893 10643 20927
rect 12725 20893 12759 20927
rect 13093 20893 13127 20927
rect 13185 20893 13219 20927
rect 13277 20893 13311 20927
rect 14105 20893 14139 20927
rect 14289 20893 14323 20927
rect 14473 20893 14507 20927
rect 14565 20893 14599 20927
rect 15117 20893 15151 20927
rect 15669 20893 15703 20927
rect 16405 20893 16439 20927
rect 18613 20893 18647 20927
rect 18889 20893 18923 20927
rect 19257 20893 19291 20927
rect 19453 20893 19487 20927
rect 19717 20893 19751 20927
rect 20085 20893 20119 20927
rect 20177 20893 20211 20927
rect 20545 20893 20579 20927
rect 20821 20893 20855 20927
rect 21005 20893 21039 20927
rect 21097 20893 21131 20927
rect 21281 20893 21315 20927
rect 21465 20893 21499 20927
rect 21833 20893 21867 20927
rect 22109 20893 22143 20927
rect 22201 20893 22235 20927
rect 22385 20893 22419 20927
rect 22477 20893 22511 20927
rect 22753 20893 22787 20927
rect 23029 20893 23063 20927
rect 23305 20893 23339 20927
rect 23397 20893 23431 20927
rect 25329 20893 25363 20927
rect 1501 20825 1535 20859
rect 1869 20825 1903 20859
rect 2237 20825 2271 20859
rect 10885 20825 10919 20859
rect 13829 20825 13863 20859
rect 18797 20825 18831 20859
rect 20729 20825 20763 20859
rect 21373 20825 21407 20859
rect 23581 20825 23615 20859
rect 24869 20825 24903 20859
rect 4905 20757 4939 20791
rect 5273 20757 5307 20791
rect 7113 20757 7147 20791
rect 12541 20757 12575 20791
rect 13737 20757 13771 20791
rect 15853 20757 15887 20791
rect 16957 20757 16991 20791
rect 17601 20757 17635 20791
rect 18429 20757 18463 20791
rect 19901 20757 19935 20791
rect 20361 20757 20395 20791
rect 21557 20757 21591 20791
rect 21925 20757 21959 20791
rect 22937 20757 22971 20791
rect 25069 20757 25103 20791
rect 25237 20757 25271 20791
rect 7665 20553 7699 20587
rect 11621 20553 11655 20587
rect 13001 20553 13035 20587
rect 14749 20553 14783 20587
rect 16037 20553 16071 20587
rect 21005 20553 21039 20587
rect 22033 20553 22067 20587
rect 22201 20553 22235 20587
rect 24225 20553 24259 20587
rect 25605 20553 25639 20587
rect 26433 20553 26467 20587
rect 1961 20485 1995 20519
rect 7113 20485 7147 20519
rect 14197 20485 14231 20519
rect 15945 20485 15979 20519
rect 19533 20485 19567 20519
rect 21281 20485 21315 20519
rect 21833 20485 21867 20519
rect 26525 20485 26559 20519
rect 2697 20417 2731 20451
rect 4813 20417 4847 20451
rect 4997 20417 5031 20451
rect 7665 20417 7699 20451
rect 11713 20417 11747 20451
rect 12265 20417 12299 20451
rect 12633 20417 12667 20451
rect 13185 20417 13219 20451
rect 13277 20417 13311 20451
rect 13461 20417 13495 20451
rect 13553 20417 13587 20451
rect 13645 20417 13679 20451
rect 13737 20417 13771 20451
rect 13921 20417 13955 20451
rect 14013 20417 14047 20451
rect 14565 20417 14599 20451
rect 15301 20417 15335 20451
rect 15393 20417 15427 20451
rect 16221 20417 16255 20451
rect 16681 20417 16715 20451
rect 17049 20417 17083 20451
rect 17601 20417 17635 20451
rect 17693 20417 17727 20451
rect 18337 20417 18371 20451
rect 18797 20417 18831 20451
rect 18889 20417 18923 20451
rect 19073 20417 19107 20451
rect 19165 20417 19199 20451
rect 21097 20417 21131 20451
rect 21373 20417 21407 20451
rect 22293 20417 22327 20451
rect 24133 20417 24167 20451
rect 25789 20417 25823 20451
rect 26065 20417 26099 20451
rect 26249 20417 26283 20451
rect 4905 20349 4939 20383
rect 5365 20349 5399 20383
rect 6193 20349 6227 20383
rect 7757 20349 7791 20383
rect 11805 20349 11839 20383
rect 12357 20349 12391 20383
rect 12541 20349 12575 20383
rect 14381 20349 14415 20383
rect 16405 20349 16439 20383
rect 19257 20349 19291 20383
rect 22569 20349 22603 20383
rect 11897 20281 11931 20315
rect 17049 20281 17083 20315
rect 18613 20213 18647 20247
rect 21097 20213 21131 20247
rect 22017 20213 22051 20247
rect 24041 20213 24075 20247
rect 4353 20009 4387 20043
rect 13093 20009 13127 20043
rect 14565 20009 14599 20043
rect 15209 20009 15243 20043
rect 15485 20009 15519 20043
rect 16589 20009 16623 20043
rect 18245 20009 18279 20043
rect 22477 20009 22511 20043
rect 23673 20009 23707 20043
rect 23857 20009 23891 20043
rect 27353 20009 27387 20043
rect 12449 19941 12483 19975
rect 20177 19941 20211 19975
rect 2145 19873 2179 19907
rect 7665 19873 7699 19907
rect 10701 19873 10735 19907
rect 10977 19873 11011 19907
rect 12541 19873 12575 19907
rect 12725 19873 12759 19907
rect 13001 19873 13035 19907
rect 15209 19873 15243 19907
rect 19073 19873 19107 19907
rect 20361 19873 20395 19907
rect 22661 19873 22695 19907
rect 25605 19873 25639 19907
rect 1409 19805 1443 19839
rect 2053 19805 2087 19839
rect 2237 19805 2271 19839
rect 2421 19805 2455 19839
rect 4261 19805 4295 19839
rect 7573 19805 7607 19839
rect 9045 19805 9079 19839
rect 9229 19805 9263 19839
rect 12909 19805 12943 19839
rect 13185 19805 13219 19839
rect 13369 19805 13403 19839
rect 13553 19805 13587 19839
rect 13645 19805 13679 19839
rect 13829 19805 13863 19839
rect 14381 19805 14415 19839
rect 14565 19805 14599 19839
rect 15117 19805 15151 19839
rect 16313 19805 16347 19839
rect 16405 19805 16439 19839
rect 18613 19805 18647 19839
rect 18705 19805 18739 19839
rect 18797 19805 18831 19839
rect 19625 19805 19659 19839
rect 19717 19805 19751 19839
rect 20085 19805 20119 19839
rect 20545 19805 20579 19839
rect 21557 19805 21591 19839
rect 21649 19805 21683 19839
rect 21925 19805 21959 19839
rect 22017 19805 22051 19839
rect 22293 19805 22327 19839
rect 22477 19805 22511 19839
rect 22753 19805 22787 19839
rect 23121 19805 23155 19839
rect 1685 19737 1719 19771
rect 3433 19737 3467 19771
rect 12817 19737 12851 19771
rect 16589 19737 16623 19771
rect 17969 19737 18003 19771
rect 18915 19737 18949 19771
rect 21833 19737 21867 19771
rect 23581 19737 23615 19771
rect 23836 19737 23870 19771
rect 24041 19737 24075 19771
rect 25881 19737 25915 19771
rect 7941 19669 7975 19703
rect 10057 19669 10091 19703
rect 13645 19669 13679 19703
rect 18429 19669 18463 19703
rect 22201 19669 22235 19703
rect 1593 19465 1627 19499
rect 3893 19465 3927 19499
rect 5365 19465 5399 19499
rect 18521 19465 18555 19499
rect 23482 19465 23516 19499
rect 27629 19465 27663 19499
rect 19349 19397 19383 19431
rect 1409 19329 1443 19363
rect 2145 19329 2179 19363
rect 2881 19329 2915 19363
rect 3065 19329 3099 19363
rect 4445 19329 4479 19363
rect 4721 19329 4755 19363
rect 5181 19329 5215 19363
rect 5365 19329 5399 19363
rect 7849 19329 7883 19363
rect 8125 19329 8159 19363
rect 8217 19329 8251 19363
rect 8677 19329 8711 19363
rect 13369 19329 13403 19363
rect 18429 19329 18463 19363
rect 18705 19329 18739 19363
rect 19257 19329 19291 19363
rect 19533 19329 19567 19363
rect 22477 19329 22511 19363
rect 22937 19329 22971 19363
rect 23305 19329 23339 19363
rect 23397 19329 23431 19363
rect 23581 19329 23615 19363
rect 27813 19329 27847 19363
rect 2053 19261 2087 19295
rect 2697 19261 2731 19295
rect 2973 19261 3007 19295
rect 3433 19261 3467 19295
rect 3525 19261 3559 19295
rect 3617 19261 3651 19295
rect 3709 19261 3743 19295
rect 5089 19261 5123 19295
rect 8585 19261 8619 19295
rect 13461 19261 13495 19295
rect 13553 19261 13587 19295
rect 13645 19261 13679 19295
rect 7941 19125 7975 19159
rect 8401 19125 8435 19159
rect 8953 19125 8987 19159
rect 13185 19125 13219 19159
rect 18889 19125 18923 19159
rect 19717 19125 19751 19159
rect 23121 19125 23155 19159
rect 9505 18921 9539 18955
rect 13093 18921 13127 18955
rect 15117 18921 15151 18955
rect 15301 18921 15335 18955
rect 17785 18921 17819 18955
rect 27813 18921 27847 18955
rect 9137 18853 9171 18887
rect 5733 18785 5767 18819
rect 22753 18785 22787 18819
rect 3433 18717 3467 18751
rect 3617 18717 3651 18751
rect 4537 18717 4571 18751
rect 4629 18717 4663 18751
rect 5273 18717 5307 18751
rect 5549 18717 5583 18751
rect 5917 18717 5951 18751
rect 6469 18717 6503 18751
rect 8217 18717 8251 18751
rect 8493 18717 8527 18751
rect 8953 18717 8987 18751
rect 9137 18717 9171 18751
rect 9413 18717 9447 18751
rect 9597 18717 9631 18751
rect 9689 18717 9723 18751
rect 9965 18717 9999 18751
rect 10149 18717 10183 18751
rect 12909 18717 12943 18751
rect 13093 18717 13127 18751
rect 14473 18717 14507 18751
rect 14657 18717 14691 18751
rect 14749 18717 14783 18751
rect 14841 18717 14875 18751
rect 15209 18717 15243 18751
rect 15761 18717 15795 18751
rect 15945 18717 15979 18751
rect 26065 18717 26099 18751
rect 8401 18649 8435 18683
rect 19073 18649 19107 18683
rect 21005 18649 21039 18683
rect 26341 18649 26375 18683
rect 3525 18581 3559 18615
rect 8315 18581 8349 18615
rect 9781 18581 9815 18615
rect 10057 18581 10091 18615
rect 13277 18581 13311 18615
rect 15853 18581 15887 18615
rect 7389 18377 7423 18411
rect 13001 18377 13035 18411
rect 13185 18377 13219 18411
rect 24593 18377 24627 18411
rect 4537 18309 4571 18343
rect 10977 18309 11011 18343
rect 3525 18241 3559 18275
rect 3709 18241 3743 18275
rect 4445 18241 4479 18275
rect 4629 18241 4663 18275
rect 4997 18241 5031 18275
rect 5273 18241 5307 18275
rect 6377 18241 6411 18275
rect 6561 18241 6595 18275
rect 7389 18241 7423 18275
rect 7665 18241 7699 18275
rect 9229 18241 9263 18275
rect 10149 18241 10183 18275
rect 10609 18241 10643 18275
rect 12817 18241 12851 18275
rect 13277 18241 13311 18275
rect 13553 18241 13587 18275
rect 14841 18241 14875 18275
rect 15301 18241 15335 18275
rect 15669 18241 15703 18275
rect 15853 18241 15887 18275
rect 16037 18241 16071 18275
rect 16313 18241 16347 18275
rect 17785 18241 17819 18275
rect 22845 18241 22879 18275
rect 4077 18173 4111 18207
rect 5825 18173 5859 18207
rect 6469 18173 6503 18207
rect 6837 18173 6871 18207
rect 7481 18173 7515 18207
rect 9137 18173 9171 18207
rect 9321 18173 9355 18207
rect 9413 18173 9447 18207
rect 12909 18173 12943 18207
rect 13461 18173 13495 18207
rect 15485 18173 15519 18207
rect 15577 18173 15611 18207
rect 23121 18173 23155 18207
rect 13921 18105 13955 18139
rect 16129 18105 16163 18139
rect 16221 18105 16255 18139
rect 7757 18037 7791 18071
rect 9597 18037 9631 18071
rect 12633 18037 12667 18071
rect 14933 18037 14967 18071
rect 15117 18037 15151 18071
rect 16497 18037 16531 18071
rect 2237 17833 2271 17867
rect 10977 17833 11011 17867
rect 13277 17833 13311 17867
rect 16773 17833 16807 17867
rect 20729 17833 20763 17867
rect 26169 17833 26203 17867
rect 8953 17765 8987 17799
rect 12449 17765 12483 17799
rect 14841 17765 14875 17799
rect 22661 17765 22695 17799
rect 9321 17697 9355 17731
rect 12633 17697 12667 17731
rect 14657 17697 14691 17731
rect 17509 17697 17543 17731
rect 18153 17697 18187 17731
rect 20361 17697 20395 17731
rect 20545 17697 20579 17731
rect 21189 17697 21223 17731
rect 22937 17697 22971 17731
rect 23397 17697 23431 17731
rect 24133 17697 24167 17731
rect 26433 17697 26467 17731
rect 2329 17629 2363 17663
rect 7665 17629 7699 17663
rect 7757 17629 7791 17663
rect 9413 17629 9447 17663
rect 9873 17629 9907 17663
rect 10241 17629 10275 17663
rect 10609 17629 10643 17663
rect 10977 17629 11011 17663
rect 11253 17629 11287 17663
rect 12725 17629 12759 17663
rect 13369 17629 13403 17663
rect 13461 17629 13495 17663
rect 13645 17629 13679 17663
rect 14933 17629 14967 17663
rect 15025 17629 15059 17663
rect 17049 17629 17083 17663
rect 17141 17629 17175 17663
rect 17877 17629 17911 17663
rect 18061 17629 18095 17663
rect 18337 17629 18371 17663
rect 18613 17629 18647 17663
rect 18889 17629 18923 17663
rect 20821 17629 20855 17663
rect 21281 17629 21315 17663
rect 22477 17629 22511 17663
rect 22569 17629 22603 17663
rect 23029 17629 23063 17663
rect 23673 17629 23707 17663
rect 23949 17629 23983 17663
rect 24225 17629 24259 17663
rect 24409 17629 24443 17663
rect 24593 17629 24627 17663
rect 8585 17561 8619 17595
rect 13001 17561 13035 17595
rect 13093 17561 13127 17595
rect 15301 17561 15335 17595
rect 17233 17561 17267 17595
rect 17351 17561 17385 17595
rect 20453 17561 20487 17595
rect 11161 17493 11195 17527
rect 13553 17493 13587 17527
rect 14933 17493 14967 17527
rect 16865 17493 16899 17527
rect 17969 17493 18003 17527
rect 18521 17493 18555 17527
rect 18797 17493 18831 17527
rect 20269 17493 20303 17527
rect 20913 17493 20947 17527
rect 24501 17493 24535 17527
rect 24685 17493 24719 17527
rect 16405 17289 16439 17323
rect 16773 17289 16807 17323
rect 19901 17289 19935 17323
rect 20545 17289 20579 17323
rect 21925 17289 21959 17323
rect 23949 17289 23983 17323
rect 1869 17221 1903 17255
rect 3065 17221 3099 17255
rect 17969 17221 18003 17255
rect 20085 17221 20119 17255
rect 24041 17221 24075 17255
rect 24409 17221 24443 17255
rect 1501 17153 1535 17187
rect 3157 17153 3191 17187
rect 3341 17153 3375 17187
rect 3801 17153 3835 17187
rect 3985 17153 4019 17187
rect 7297 17153 7331 17187
rect 8033 17153 8067 17187
rect 8585 17153 8619 17187
rect 9873 17153 9907 17187
rect 10057 17153 10091 17187
rect 11805 17153 11839 17187
rect 11897 17153 11931 17187
rect 11989 17153 12023 17187
rect 12173 17153 12207 17187
rect 14565 17153 14599 17187
rect 14749 17153 14783 17187
rect 15761 17153 15795 17187
rect 15945 17153 15979 17187
rect 16129 17153 16163 17187
rect 16221 17153 16255 17187
rect 16497 17153 16531 17187
rect 16681 17153 16715 17187
rect 16957 17153 16991 17187
rect 17233 17153 17267 17187
rect 17693 17153 17727 17187
rect 19717 17153 19751 17187
rect 19993 17153 20027 17187
rect 20269 17153 20303 17187
rect 20361 17153 20395 17187
rect 20637 17153 20671 17187
rect 20821 17153 20855 17187
rect 20913 17153 20947 17187
rect 21005 17153 21039 17187
rect 21557 17153 21591 17187
rect 21833 17153 21867 17187
rect 22017 17153 22051 17187
rect 23213 17153 23247 17187
rect 23397 17153 23431 17187
rect 23489 17153 23523 17187
rect 23765 17153 23799 17187
rect 24225 17153 24259 17187
rect 24685 17153 24719 17187
rect 24777 17153 24811 17187
rect 2237 17085 2271 17119
rect 6377 17085 6411 17119
rect 7389 17085 7423 17119
rect 10885 17085 10919 17119
rect 12265 17085 12299 17119
rect 12541 17085 12575 17119
rect 15025 17085 15059 17119
rect 15301 17085 15335 17119
rect 17049 17085 17083 17119
rect 21281 17085 21315 17119
rect 23581 17085 23615 17119
rect 6837 17017 6871 17051
rect 11713 17017 11747 17051
rect 14933 17017 14967 17051
rect 16221 17017 16255 17051
rect 21189 17017 21223 17051
rect 24501 17017 24535 17051
rect 3341 16949 3375 16983
rect 3893 16949 3927 16983
rect 9505 16949 9539 16983
rect 14013 16949 14047 16983
rect 14841 16949 14875 16983
rect 15393 16949 15427 16983
rect 15669 16949 15703 16983
rect 15853 16949 15887 16983
rect 16957 16949 16991 16983
rect 17417 16949 17451 16983
rect 20085 16949 20119 16983
rect 21373 16949 21407 16983
rect 21465 16949 21499 16983
rect 2421 16745 2455 16779
rect 7757 16745 7791 16779
rect 9321 16745 9355 16779
rect 13461 16745 13495 16779
rect 17417 16745 17451 16779
rect 17739 16745 17773 16779
rect 18153 16745 18187 16779
rect 26341 16745 26375 16779
rect 1961 16609 1995 16643
rect 2237 16609 2271 16643
rect 3157 16609 3191 16643
rect 3249 16609 3283 16643
rect 3433 16609 3467 16643
rect 4077 16609 4111 16643
rect 13001 16609 13035 16643
rect 13093 16609 13127 16643
rect 17233 16609 17267 16643
rect 17877 16609 17911 16643
rect 20545 16609 20579 16643
rect 20729 16609 20763 16643
rect 25881 16609 25915 16643
rect 26157 16609 26191 16643
rect 1869 16541 1903 16575
rect 2329 16531 2363 16565
rect 2513 16541 2547 16575
rect 2973 16541 3007 16575
rect 3065 16541 3099 16575
rect 4169 16541 4203 16575
rect 5089 16541 5123 16575
rect 5273 16541 5307 16575
rect 5457 16541 5491 16575
rect 6009 16541 6043 16575
rect 8033 16541 8067 16575
rect 8585 16541 8619 16575
rect 9137 16541 9171 16575
rect 9321 16541 9355 16575
rect 12081 16541 12115 16575
rect 12265 16541 12299 16575
rect 12449 16541 12483 16575
rect 12725 16541 12759 16575
rect 12909 16541 12943 16575
rect 13277 16541 13311 16575
rect 17509 16541 17543 16575
rect 17601 16541 17635 16575
rect 18061 16541 18095 16575
rect 18337 16541 18371 16575
rect 18521 16541 18555 16575
rect 18613 16541 18647 16575
rect 18705 16541 18739 16575
rect 18889 16541 18923 16575
rect 20453 16541 20487 16575
rect 21005 16541 21039 16575
rect 21281 16541 21315 16575
rect 21373 16541 21407 16575
rect 21557 16541 21591 16575
rect 22109 16541 22143 16575
rect 22201 16541 22235 16575
rect 23489 16541 23523 16575
rect 7757 16473 7791 16507
rect 8401 16473 8435 16507
rect 12357 16473 12391 16507
rect 20729 16473 20763 16507
rect 21189 16473 21223 16507
rect 26617 16473 26651 16507
rect 4905 16405 4939 16439
rect 5181 16405 5215 16439
rect 7941 16405 7975 16439
rect 8769 16405 8803 16439
rect 12633 16405 12667 16439
rect 17233 16405 17267 16439
rect 18061 16405 18095 16439
rect 20821 16405 20855 16439
rect 21373 16405 21407 16439
rect 23397 16405 23431 16439
rect 24409 16405 24443 16439
rect 17693 16201 17727 16235
rect 22477 16201 22511 16235
rect 23489 16201 23523 16235
rect 25329 16201 25363 16235
rect 8677 16133 8711 16167
rect 12817 16133 12851 16167
rect 18153 16133 18187 16167
rect 23765 16133 23799 16167
rect 25605 16133 25639 16167
rect 1869 16065 1903 16099
rect 3893 16065 3927 16099
rect 4629 16065 4663 16099
rect 4905 16065 4939 16099
rect 5365 16065 5399 16099
rect 6745 16065 6779 16099
rect 7481 16065 7515 16099
rect 9045 16065 9079 16099
rect 9781 16065 9815 16099
rect 9965 16065 9999 16099
rect 13093 16065 13127 16099
rect 17877 16065 17911 16099
rect 18521 16065 18555 16099
rect 20545 16065 20579 16099
rect 20821 16065 20855 16099
rect 21281 16065 21315 16099
rect 21465 16065 21499 16099
rect 22661 16065 22695 16099
rect 22753 16065 22787 16099
rect 22937 16065 22971 16099
rect 23029 16065 23063 16099
rect 23305 16065 23339 16099
rect 23581 16065 23615 16099
rect 23673 16065 23707 16099
rect 23949 16065 23983 16099
rect 1961 15997 1995 16031
rect 4537 15997 4571 16031
rect 8861 15997 8895 16031
rect 13001 15997 13035 16031
rect 17969 15997 18003 16031
rect 18245 15997 18279 16031
rect 21097 15997 21131 16031
rect 23121 15997 23155 16031
rect 9045 15929 9079 15963
rect 13277 15929 13311 15963
rect 18429 15929 18463 15963
rect 2145 15861 2179 15895
rect 8217 15861 8251 15895
rect 12817 15861 12851 15895
rect 18153 15861 18187 15895
rect 18521 15861 18555 15895
rect 19257 15861 19291 15895
rect 20637 15861 20671 15895
rect 21005 15861 21039 15895
rect 21281 15861 21315 15895
rect 24133 15861 24167 15895
rect 7573 15657 7607 15691
rect 20913 15657 20947 15691
rect 21097 15657 21131 15691
rect 23489 15657 23523 15691
rect 23949 15657 23983 15691
rect 24409 15657 24443 15691
rect 24593 15657 24627 15691
rect 8677 15589 8711 15623
rect 19441 15589 19475 15623
rect 20361 15589 20395 15623
rect 21373 15589 21407 15623
rect 23121 15589 23155 15623
rect 23857 15589 23891 15623
rect 24869 15589 24903 15623
rect 4537 15521 4571 15555
rect 8033 15521 8067 15555
rect 19625 15521 19659 15555
rect 1409 15453 1443 15487
rect 2789 15453 2823 15487
rect 3065 15453 3099 15487
rect 4445 15453 4479 15487
rect 4905 15453 4939 15487
rect 5089 15453 5123 15487
rect 7757 15453 7791 15487
rect 7849 15453 7883 15487
rect 8125 15453 8159 15487
rect 8585 15453 8619 15487
rect 8769 15453 8803 15487
rect 9321 15453 9355 15487
rect 9873 15453 9907 15487
rect 19441 15453 19475 15487
rect 19809 15453 19843 15487
rect 20545 15453 20579 15487
rect 20729 15453 20763 15487
rect 21281 15453 21315 15487
rect 21465 15453 21499 15487
rect 21557 15453 21591 15487
rect 21741 15453 21775 15487
rect 21925 15453 21959 15487
rect 22937 15453 22971 15487
rect 23765 15453 23799 15487
rect 24041 15453 24075 15487
rect 24225 15453 24259 15487
rect 25053 15453 25087 15487
rect 25145 15453 25179 15487
rect 1685 15385 1719 15419
rect 4997 15385 5031 15419
rect 21005 15385 21039 15419
rect 21833 15385 21867 15419
rect 24777 15385 24811 15419
rect 24869 15385 24903 15419
rect 3433 15317 3467 15351
rect 4813 15317 4847 15351
rect 24577 15317 24611 15351
rect 2881 15113 2915 15147
rect 12081 15113 12115 15147
rect 15117 15113 15151 15147
rect 18889 15113 18923 15147
rect 20821 15113 20855 15147
rect 9873 15045 9907 15079
rect 11805 15045 11839 15079
rect 15301 15045 15335 15079
rect 2789 14977 2823 15011
rect 2973 14977 3007 15011
rect 3249 14977 3283 15011
rect 8217 14977 8251 15011
rect 8401 14977 8435 15011
rect 11529 14977 11563 15011
rect 11713 14977 11747 15011
rect 11897 14977 11931 15011
rect 12633 14977 12667 15011
rect 13001 14977 13035 15011
rect 18429 14977 18463 15011
rect 18705 14977 18739 15011
rect 21189 14977 21223 15011
rect 24317 14977 24351 15011
rect 5457 14909 5491 14943
rect 12173 14909 12207 14943
rect 12725 14909 12759 14943
rect 12909 14909 12943 14943
rect 15209 14909 15243 14943
rect 15393 14909 15427 14943
rect 15669 14909 15703 14943
rect 18521 14909 18555 14943
rect 21097 14909 21131 14943
rect 5733 14841 5767 14875
rect 12265 14841 12299 14875
rect 3341 14773 3375 14807
rect 5917 14773 5951 14807
rect 15577 14773 15611 14807
rect 18705 14773 18739 14807
rect 24225 14773 24259 14807
rect 13093 14569 13127 14603
rect 15577 14569 15611 14603
rect 27629 14569 27663 14603
rect 3985 14501 4019 14535
rect 6469 14501 6503 14535
rect 14703 14501 14737 14535
rect 15761 14501 15795 14535
rect 16957 14501 16991 14535
rect 25329 14501 25363 14535
rect 3525 14433 3559 14467
rect 4077 14433 4111 14467
rect 4353 14433 4387 14467
rect 6101 14433 6135 14467
rect 7021 14433 7055 14467
rect 11069 14433 11103 14467
rect 13829 14433 13863 14467
rect 15209 14433 15243 14467
rect 17049 14433 17083 14467
rect 17141 14433 17175 14467
rect 24501 14433 24535 14467
rect 2789 14365 2823 14399
rect 3249 14365 3283 14399
rect 3893 14365 3927 14399
rect 4169 14365 4203 14399
rect 5089 14365 5123 14399
rect 5457 14365 5491 14399
rect 6193 14365 6227 14399
rect 6745 14365 6779 14399
rect 11161 14365 11195 14399
rect 11253 14365 11287 14399
rect 13277 14365 13311 14399
rect 13369 14365 13403 14399
rect 13553 14365 13587 14399
rect 13645 14365 13679 14399
rect 13737 14365 13771 14399
rect 14289 14365 14323 14399
rect 14473 14365 14507 14399
rect 14565 14365 14599 14399
rect 14841 14365 14875 14399
rect 15025 14365 15059 14399
rect 15117 14365 15151 14399
rect 15393 14365 15427 14399
rect 16681 14365 16715 14399
rect 16773 14365 16807 14399
rect 16957 14365 16991 14399
rect 20361 14365 20395 14399
rect 24593 14365 24627 14399
rect 27813 14365 27847 14399
rect 11529 14297 11563 14331
rect 14933 14297 14967 14331
rect 16037 14297 16071 14331
rect 23305 14297 23339 14331
rect 25145 14297 25179 14331
rect 13001 14229 13035 14263
rect 14381 14229 14415 14263
rect 20269 14229 20303 14263
rect 23581 14229 23615 14263
rect 24961 14229 24995 14263
rect 2789 14025 2823 14059
rect 3617 14025 3651 14059
rect 17417 14025 17451 14059
rect 19257 14025 19291 14059
rect 25697 14025 25731 14059
rect 1685 13957 1719 13991
rect 11805 13957 11839 13991
rect 13461 13957 13495 13991
rect 14657 13957 14691 13991
rect 17049 13957 17083 13991
rect 18061 13957 18095 13991
rect 19993 13957 20027 13991
rect 21097 13957 21131 13991
rect 21465 13957 21499 13991
rect 22753 13957 22787 13991
rect 1409 13889 1443 13923
rect 2237 13889 2271 13923
rect 3065 13889 3099 13923
rect 3157 13889 3191 13923
rect 3433 13889 3467 13923
rect 3617 13889 3651 13923
rect 3709 13889 3743 13923
rect 3893 13889 3927 13923
rect 4169 13889 4203 13923
rect 4353 13889 4387 13923
rect 5825 13889 5859 13923
rect 6929 13889 6963 13923
rect 7205 13889 7239 13923
rect 7573 13889 7607 13923
rect 9413 13889 9447 13923
rect 9597 13889 9631 13923
rect 9689 13889 9723 13923
rect 11529 13889 11563 13923
rect 13737 13889 13771 13923
rect 14197 13889 14231 13923
rect 14381 13889 14415 13923
rect 16865 13889 16899 13923
rect 17141 13889 17175 13923
rect 17233 13889 17267 13923
rect 18613 13889 18647 13923
rect 18705 13889 18739 13923
rect 18981 13889 19015 13923
rect 19073 13889 19107 13923
rect 19533 13889 19567 13923
rect 19809 13889 19843 13923
rect 20085 13889 20119 13923
rect 20350 13889 20384 13923
rect 20729 13889 20763 13923
rect 20913 13889 20947 13923
rect 21189 13889 21223 13923
rect 21649 13889 21683 13923
rect 22201 13889 22235 13923
rect 22293 13889 22327 13923
rect 22477 13889 22511 13923
rect 22569 13889 22603 13923
rect 22845 13889 22879 13923
rect 23029 13889 23063 13923
rect 23397 13889 23431 13923
rect 23949 13889 23983 13923
rect 2329 13821 2363 13855
rect 2605 13821 2639 13855
rect 2973 13821 3007 13855
rect 3249 13821 3283 13855
rect 3801 13821 3835 13855
rect 5917 13821 5951 13855
rect 8677 13821 8711 13855
rect 18245 13821 18279 13855
rect 18337 13821 18371 13855
rect 18429 13821 18463 13855
rect 19441 13821 19475 13855
rect 20545 13821 20579 13855
rect 20637 13821 20671 13855
rect 21281 13821 21315 13855
rect 23581 13821 23615 13855
rect 23857 13821 23891 13855
rect 24225 13821 24259 13855
rect 6193 13753 6227 13787
rect 7481 13753 7515 13787
rect 8953 13753 8987 13787
rect 14013 13753 14047 13787
rect 18153 13753 18187 13787
rect 18797 13753 18831 13787
rect 23765 13753 23799 13787
rect 4353 13685 4387 13719
rect 9137 13685 9171 13719
rect 9229 13685 9263 13719
rect 13277 13685 13311 13719
rect 13829 13685 13863 13719
rect 13921 13685 13955 13719
rect 16129 13685 16163 13719
rect 19625 13685 19659 13719
rect 20177 13685 20211 13719
rect 8769 13481 8803 13515
rect 10241 13481 10275 13515
rect 13001 13481 13035 13515
rect 14933 13481 14967 13515
rect 15485 13481 15519 13515
rect 18521 13481 18555 13515
rect 21465 13481 21499 13515
rect 21557 13481 21591 13515
rect 22385 13481 22419 13515
rect 24409 13481 24443 13515
rect 6929 13413 6963 13447
rect 13185 13413 13219 13447
rect 18613 13413 18647 13447
rect 24777 13413 24811 13447
rect 2973 13345 3007 13379
rect 4721 13345 4755 13379
rect 9137 13345 9171 13379
rect 12081 13345 12115 13379
rect 15853 13345 15887 13379
rect 15945 13345 15979 13379
rect 16681 13345 16715 13379
rect 18705 13345 18739 13379
rect 21925 13345 21959 13379
rect 22937 13345 22971 13379
rect 23213 13345 23247 13379
rect 2881 13277 2915 13311
rect 3341 13277 3375 13311
rect 3525 13277 3559 13311
rect 4629 13277 4663 13311
rect 6929 13277 6963 13311
rect 7205 13277 7239 13311
rect 8217 13277 8251 13311
rect 8309 13277 8343 13311
rect 8493 13277 8527 13311
rect 8585 13277 8619 13311
rect 9229 13277 9263 13311
rect 10149 13277 10183 13311
rect 11989 13277 12023 13311
rect 12725 13277 12759 13311
rect 12817 13277 12851 13311
rect 13001 13277 13035 13311
rect 13093 13277 13127 13311
rect 13277 13277 13311 13311
rect 13553 13277 13587 13311
rect 14657 13277 14691 13311
rect 14841 13277 14875 13311
rect 15117 13277 15151 13311
rect 15301 13277 15335 13311
rect 15393 13277 15427 13311
rect 15669 13277 15703 13311
rect 16037 13277 16071 13311
rect 16221 13277 16255 13311
rect 18429 13277 18463 13311
rect 19441 13277 19475 13311
rect 19625 13277 19659 13311
rect 19717 13277 19751 13311
rect 21557 13277 21591 13311
rect 21741 13277 21775 13311
rect 22017 13277 22051 13311
rect 22109 13277 22143 13311
rect 22201 13277 22235 13311
rect 22845 13277 22879 13311
rect 24593 13277 24627 13311
rect 24685 13277 24719 13311
rect 24869 13277 24903 13311
rect 3433 13209 3467 13243
rect 7113 13209 7147 13243
rect 11621 13209 11655 13243
rect 11713 13209 11747 13243
rect 14749 13209 14783 13243
rect 16313 13209 16347 13243
rect 16497 13209 16531 13243
rect 19533 13209 19567 13243
rect 19993 13209 20027 13243
rect 3249 13141 3283 13175
rect 5273 13141 5307 13175
rect 10057 13141 10091 13175
rect 12265 13141 12299 13175
rect 13737 13141 13771 13175
rect 2237 12937 2271 12971
rect 6561 12937 6595 12971
rect 7297 12937 7331 12971
rect 13201 12937 13235 12971
rect 13369 12937 13403 12971
rect 15761 12937 15795 12971
rect 18705 12937 18739 12971
rect 22201 12937 22235 12971
rect 13001 12869 13035 12903
rect 20085 12869 20119 12903
rect 22937 12869 22971 12903
rect 24133 12869 24167 12903
rect 2237 12801 2271 12835
rect 2421 12801 2455 12835
rect 5181 12801 5215 12835
rect 6377 12801 6411 12835
rect 6561 12801 6595 12835
rect 7205 12801 7239 12835
rect 7389 12801 7423 12835
rect 8585 12801 8619 12835
rect 9413 12801 9447 12835
rect 15117 12801 15151 12835
rect 15393 12801 15427 12835
rect 15577 12801 15611 12835
rect 16037 12801 16071 12835
rect 17325 12801 17359 12835
rect 18797 12801 18831 12835
rect 19717 12801 19751 12835
rect 20361 12801 20395 12835
rect 20729 12801 20763 12835
rect 20913 12801 20947 12835
rect 21005 12801 21039 12835
rect 21189 12801 21223 12835
rect 21833 12801 21867 12835
rect 22017 12801 22051 12835
rect 22477 12801 22511 12835
rect 23397 12801 23431 12835
rect 23857 12801 23891 12835
rect 24225 12801 24259 12835
rect 6193 12733 6227 12767
rect 7757 12733 7791 12767
rect 9505 12733 9539 12767
rect 10057 12733 10091 12767
rect 22293 12733 22327 12767
rect 23305 12733 23339 12767
rect 23673 12733 23707 12767
rect 16221 12665 16255 12699
rect 22661 12665 22695 12699
rect 13185 12597 13219 12631
rect 15209 12597 15243 12631
rect 17049 12597 17083 12631
rect 20085 12597 20119 12631
rect 20269 12597 20303 12631
rect 20729 12597 20763 12631
rect 21097 12597 21131 12631
rect 23213 12597 23247 12631
rect 23581 12597 23615 12631
rect 12357 12393 12391 12427
rect 15577 12393 15611 12427
rect 15853 12393 15887 12427
rect 19257 12393 19291 12427
rect 15761 12325 15795 12359
rect 19625 12325 19659 12359
rect 1961 12257 1995 12291
rect 2237 12257 2271 12291
rect 2421 12257 2455 12291
rect 6561 12257 6595 12291
rect 7481 12257 7515 12291
rect 12725 12257 12759 12291
rect 16037 12257 16071 12291
rect 19533 12257 19567 12291
rect 1869 12189 1903 12223
rect 2513 12189 2547 12223
rect 6107 12189 6141 12223
rect 6285 12189 6319 12223
rect 6653 12189 6687 12223
rect 12541 12189 12575 12223
rect 12633 12189 12667 12223
rect 12817 12189 12851 12223
rect 16129 12189 16163 12223
rect 17049 12189 17083 12223
rect 18797 12189 18831 12223
rect 19441 12189 19475 12223
rect 19717 12189 19751 12223
rect 19901 12189 19935 12223
rect 15393 12121 15427 12155
rect 15593 12121 15627 12155
rect 15853 12121 15887 12155
rect 16773 12121 16807 12155
rect 20269 12121 20303 12155
rect 2881 12053 2915 12087
rect 6285 12053 6319 12087
rect 16313 12053 16347 12087
rect 16497 12053 16531 12087
rect 21557 12053 21591 12087
rect 9597 11849 9631 11883
rect 12541 11849 12575 11883
rect 13185 11849 13219 11883
rect 15577 11849 15611 11883
rect 19993 11849 20027 11883
rect 23673 11849 23707 11883
rect 25421 11849 25455 11883
rect 4721 11781 4755 11815
rect 8953 11781 8987 11815
rect 10977 11781 11011 11815
rect 11177 11781 11211 11815
rect 14013 11781 14047 11815
rect 14105 11781 14139 11815
rect 16037 11781 16071 11815
rect 18613 11781 18647 11815
rect 19073 11781 19107 11815
rect 23949 11781 23983 11815
rect 1409 11713 1443 11747
rect 3893 11713 3927 11747
rect 4353 11723 4387 11757
rect 4537 11713 4571 11747
rect 4629 11713 4663 11747
rect 4905 11713 4939 11747
rect 5181 11713 5215 11747
rect 5365 11713 5399 11747
rect 8493 11713 8527 11747
rect 8677 11713 8711 11747
rect 8769 11713 8803 11747
rect 9137 11713 9171 11747
rect 9413 11713 9447 11747
rect 9597 11713 9631 11747
rect 9689 11713 9723 11747
rect 9873 11713 9907 11747
rect 12725 11713 12759 11747
rect 12817 11713 12851 11747
rect 13001 11713 13035 11747
rect 13093 11713 13127 11747
rect 13369 11713 13403 11747
rect 13553 11713 13587 11747
rect 13645 11713 13679 11747
rect 13829 11713 13863 11747
rect 14197 11713 14231 11747
rect 14657 11713 14691 11747
rect 15301 11713 15335 11747
rect 15393 11713 15427 11747
rect 15669 11713 15703 11747
rect 15945 11713 15979 11747
rect 16129 11713 16163 11747
rect 16313 11713 16347 11747
rect 16405 11713 16439 11747
rect 17049 11713 17083 11747
rect 18061 11713 18095 11747
rect 18153 11713 18187 11747
rect 18337 11713 18371 11747
rect 18429 11713 18463 11747
rect 19533 11713 19567 11747
rect 20545 11713 20579 11747
rect 23857 11713 23891 11747
rect 24041 11713 24075 11747
rect 24225 11713 24259 11747
rect 24317 11713 24351 11747
rect 24593 11713 24627 11747
rect 25697 11713 25731 11747
rect 1685 11645 1719 11679
rect 3801 11645 3835 11679
rect 4445 11645 4479 11679
rect 8585 11645 8619 11679
rect 15485 11645 15519 11679
rect 19625 11645 19659 11679
rect 20269 11645 20303 11679
rect 4261 11577 4295 11611
rect 11345 11577 11379 11611
rect 19901 11577 19935 11611
rect 9873 11509 9907 11543
rect 11161 11509 11195 11543
rect 14381 11509 14415 11543
rect 14749 11509 14783 11543
rect 15761 11509 15795 11543
rect 18797 11509 18831 11543
rect 20177 11509 20211 11543
rect 24501 11509 24535 11543
rect 4353 11305 4387 11339
rect 10333 11305 10367 11339
rect 12173 11305 12207 11339
rect 12725 11305 12759 11339
rect 13185 11305 13219 11339
rect 15577 11305 15611 11339
rect 19809 11305 19843 11339
rect 23489 11305 23523 11339
rect 24225 11305 24259 11339
rect 24666 11305 24700 11339
rect 26157 11305 26191 11339
rect 5457 11237 5491 11271
rect 7205 11237 7239 11271
rect 23857 11237 23891 11271
rect 3065 11169 3099 11203
rect 3893 11169 3927 11203
rect 3985 11169 4019 11203
rect 4905 11169 4939 11203
rect 7573 11169 7607 11203
rect 9321 11169 9355 11203
rect 13093 11169 13127 11203
rect 16589 11169 16623 11203
rect 18705 11169 18739 11203
rect 19533 11169 19567 11203
rect 21557 11169 21591 11203
rect 24409 11169 24443 11203
rect 2973 11101 3007 11135
rect 3157 11101 3191 11135
rect 4077 11101 4111 11135
rect 4169 11101 4203 11135
rect 4997 11101 5031 11135
rect 5457 11101 5491 11135
rect 5641 11101 5675 11135
rect 7481 11101 7515 11135
rect 9505 11101 9539 11135
rect 9689 11101 9723 11135
rect 10609 11101 10643 11135
rect 11805 11101 11839 11135
rect 11989 11101 12023 11135
rect 12081 11101 12115 11135
rect 12265 11101 12299 11135
rect 12909 11101 12943 11135
rect 13277 11101 13311 11135
rect 13553 11101 13587 11135
rect 13737 11101 13771 11135
rect 15393 11101 15427 11135
rect 15577 11101 15611 11135
rect 15669 11101 15703 11135
rect 15853 11101 15887 11135
rect 15945 11101 15979 11135
rect 16037 11101 16071 11135
rect 16313 11101 16347 11135
rect 18337 11101 18371 11135
rect 19349 11101 19383 11135
rect 19441 11101 19475 11135
rect 19625 11101 19659 11135
rect 21097 11101 21131 11135
rect 21281 11101 21315 11135
rect 21373 11101 21407 11135
rect 21649 11101 21683 11135
rect 23213 11101 23247 11135
rect 23581 11101 23615 11135
rect 23765 11101 23799 11135
rect 23949 11101 23983 11135
rect 24041 11101 24075 11135
rect 6929 11033 6963 11067
rect 9873 11033 9907 11067
rect 10517 11033 10551 11067
rect 10701 11033 10735 11067
rect 10885 11033 10919 11067
rect 11897 11033 11931 11067
rect 13185 11033 13219 11067
rect 13645 11033 13679 11067
rect 18521 11033 18555 11067
rect 23305 11033 23339 11067
rect 23489 11033 23523 11067
rect 5365 10965 5399 10999
rect 9597 10965 9631 10999
rect 12449 10965 12483 10999
rect 13369 10965 13403 10999
rect 16221 10965 16255 10999
rect 18061 10965 18095 10999
rect 20913 10965 20947 10999
rect 3249 10761 3283 10795
rect 5825 10761 5859 10795
rect 8677 10761 8711 10795
rect 15485 10761 15519 10795
rect 16405 10761 16439 10795
rect 18153 10761 18187 10795
rect 24517 10761 24551 10795
rect 9689 10693 9723 10727
rect 10057 10693 10091 10727
rect 11621 10693 11655 10727
rect 16037 10693 16071 10727
rect 17417 10693 17451 10727
rect 20821 10693 20855 10727
rect 21005 10693 21039 10727
rect 23765 10693 23799 10727
rect 24317 10693 24351 10727
rect 25145 10693 25179 10727
rect 1869 10625 1903 10659
rect 2697 10625 2731 10659
rect 3157 10625 3191 10659
rect 3341 10625 3375 10659
rect 6039 10625 6073 10659
rect 6204 10625 6238 10659
rect 6561 10625 6595 10659
rect 7389 10625 7423 10659
rect 8585 10625 8619 10659
rect 8769 10625 8803 10659
rect 9229 10625 9263 10659
rect 9413 10625 9447 10659
rect 9505 10625 9539 10659
rect 9873 10625 9907 10659
rect 9965 10625 9999 10659
rect 10149 10625 10183 10659
rect 11529 10625 11563 10659
rect 11713 10625 11747 10659
rect 11805 10625 11839 10659
rect 11897 10625 11931 10659
rect 12081 10625 12115 10659
rect 12173 10625 12207 10659
rect 12357 10625 12391 10659
rect 12633 10625 12667 10659
rect 12817 10625 12851 10659
rect 13001 10625 13035 10659
rect 13185 10625 13219 10659
rect 14013 10625 14047 10659
rect 14197 10625 14231 10659
rect 14473 10625 14507 10659
rect 15117 10625 15151 10659
rect 15301 10625 15335 10659
rect 16221 10625 16255 10659
rect 16497 10625 16531 10659
rect 16681 10625 16715 10659
rect 16865 10625 16899 10659
rect 17233 10625 17267 10659
rect 17509 10625 17543 10659
rect 17602 10625 17636 10659
rect 17785 10625 17819 10659
rect 17877 10625 17911 10659
rect 17974 10625 18008 10659
rect 20177 10625 20211 10659
rect 20453 10625 20487 10659
rect 20637 10625 20671 10659
rect 20913 10625 20947 10659
rect 21189 10625 21223 10659
rect 21281 10625 21315 10659
rect 21465 10625 21499 10659
rect 21557 10625 21591 10659
rect 24041 10625 24075 10659
rect 24777 10625 24811 10659
rect 24961 10625 24995 10659
rect 1961 10557 1995 10591
rect 2605 10557 2639 10591
rect 6469 10557 6503 10591
rect 7481 10557 7515 10591
rect 9045 10557 9079 10591
rect 12909 10557 12943 10591
rect 13369 10557 13403 10591
rect 16951 10557 16985 10591
rect 17049 10557 17083 10591
rect 23857 10557 23891 10591
rect 2237 10489 2271 10523
rect 6929 10489 6963 10523
rect 7757 10489 7791 10523
rect 14657 10489 14691 10523
rect 24225 10489 24259 10523
rect 3065 10421 3099 10455
rect 15117 10421 15151 10455
rect 20269 10421 20303 10455
rect 23857 10421 23891 10455
rect 24501 10421 24535 10455
rect 24685 10421 24719 10455
rect 7757 10217 7791 10251
rect 8493 10217 8527 10251
rect 12173 10217 12207 10251
rect 13001 10217 13035 10251
rect 13185 10217 13219 10251
rect 14197 10217 14231 10251
rect 14749 10217 14783 10251
rect 16405 10217 16439 10251
rect 16957 10217 16991 10251
rect 20453 10217 20487 10251
rect 24501 10217 24535 10251
rect 24869 10217 24903 10251
rect 3157 10149 3191 10183
rect 18705 10149 18739 10183
rect 2697 10081 2731 10115
rect 4077 10081 4111 10115
rect 7941 10081 7975 10115
rect 8953 10081 8987 10115
rect 13829 10081 13863 10115
rect 16681 10081 16715 10115
rect 18429 10081 18463 10115
rect 18613 10081 18647 10115
rect 19809 10081 19843 10115
rect 20821 10081 20855 10115
rect 25053 10081 25087 10115
rect 25329 10081 25363 10115
rect 2789 10013 2823 10047
rect 3985 10013 4019 10047
rect 4445 10013 4479 10047
rect 4629 10013 4663 10047
rect 7665 10013 7699 10047
rect 7849 10013 7883 10047
rect 8125 10013 8159 10047
rect 8217 10013 8251 10047
rect 8309 9991 8343 10025
rect 8401 10013 8435 10047
rect 9321 10013 9355 10047
rect 9505 10013 9539 10047
rect 9781 10013 9815 10047
rect 11621 10013 11655 10047
rect 11805 10013 11839 10047
rect 11989 10013 12023 10047
rect 12265 10013 12299 10047
rect 12449 10013 12483 10047
rect 12725 10013 12759 10047
rect 13277 10013 13311 10047
rect 13461 10013 13495 10047
rect 13553 10013 13587 10047
rect 13737 10013 13771 10047
rect 14381 10013 14415 10047
rect 14565 10013 14599 10047
rect 16497 10013 16531 10047
rect 16773 10013 16807 10047
rect 16865 10013 16899 10047
rect 17059 10013 17093 10047
rect 18337 10013 18371 10047
rect 18797 10013 18831 10047
rect 19717 10013 19751 10047
rect 19901 10013 19935 10047
rect 20177 10013 20211 10047
rect 20545 10013 20579 10047
rect 24409 10013 24443 10047
rect 24593 10013 24627 10047
rect 24961 10013 24995 10047
rect 4537 9945 4571 9979
rect 7941 9945 7975 9979
rect 9597 9945 9631 9979
rect 9965 9945 9999 9979
rect 11897 9945 11931 9979
rect 12817 9945 12851 9979
rect 13033 9945 13067 9979
rect 14105 9945 14139 9979
rect 18705 9945 18739 9979
rect 19257 9945 19291 9979
rect 19441 9945 19475 9979
rect 19625 9945 19659 9979
rect 20453 9945 20487 9979
rect 4353 9877 4387 9911
rect 8677 9877 8711 9911
rect 9321 9877 9355 9911
rect 12633 9877 12667 9911
rect 20269 9877 20303 9911
rect 22293 9877 22327 9911
rect 26801 9877 26835 9911
rect 9137 9673 9171 9707
rect 18521 9673 18555 9707
rect 21833 9673 21867 9707
rect 8769 9605 8803 9639
rect 8985 9605 9019 9639
rect 18889 9605 18923 9639
rect 20913 9605 20947 9639
rect 21113 9605 21147 9639
rect 12173 9537 12207 9571
rect 12265 9537 12299 9571
rect 12408 9537 12442 9571
rect 12541 9537 12575 9571
rect 12909 9537 12943 9571
rect 13093 9537 13127 9571
rect 13369 9537 13403 9571
rect 13461 9537 13495 9571
rect 13645 9537 13679 9571
rect 18153 9537 18187 9571
rect 18705 9537 18739 9571
rect 18981 9537 19015 9571
rect 22109 9537 22143 9571
rect 22201 9537 22235 9571
rect 22569 9537 22603 9571
rect 24041 9537 24075 9571
rect 24225 9537 24259 9571
rect 18245 9469 18279 9503
rect 22385 9469 22419 9503
rect 13001 9401 13035 9435
rect 13461 9401 13495 9435
rect 18981 9401 19015 9435
rect 21281 9401 21315 9435
rect 22293 9401 22327 9435
rect 8953 9333 8987 9367
rect 11989 9333 12023 9367
rect 12633 9333 12667 9367
rect 13185 9333 13219 9367
rect 21097 9333 21131 9367
rect 24225 9333 24259 9367
rect 24501 9333 24535 9367
rect 6285 9129 6319 9163
rect 8217 9129 8251 9163
rect 11897 9129 11931 9163
rect 13093 9129 13127 9163
rect 16865 9129 16899 9163
rect 23397 9129 23431 9163
rect 24869 9129 24903 9163
rect 25145 9129 25179 9163
rect 17417 9061 17451 9095
rect 24961 9061 24995 9095
rect 4997 8993 5031 9027
rect 9965 8993 9999 9027
rect 24133 8993 24167 9027
rect 24777 8993 24811 9027
rect 5089 8925 5123 8959
rect 5825 8925 5859 8959
rect 5917 8925 5951 8959
rect 6009 8925 6043 8959
rect 6101 8925 6135 8959
rect 8125 8925 8159 8959
rect 8309 8925 8343 8959
rect 9689 8925 9723 8959
rect 9781 8925 9815 8959
rect 12081 8925 12115 8959
rect 12265 8925 12299 8959
rect 12357 8925 12391 8959
rect 12449 8925 12483 8959
rect 13093 8925 13127 8959
rect 13277 8925 13311 8959
rect 17141 8925 17175 8959
rect 17233 8925 17267 8959
rect 23029 8925 23063 8959
rect 23121 8925 23155 8959
rect 23581 8925 23615 8959
rect 23673 8925 23707 8959
rect 23949 8925 23983 8959
rect 24041 8925 24075 8959
rect 24225 8925 24259 8959
rect 24593 8925 24627 8959
rect 24869 8925 24903 8959
rect 16681 8857 16715 8891
rect 16881 8857 16915 8891
rect 17417 8857 17451 8891
rect 23765 8857 23799 8891
rect 25113 8857 25147 8891
rect 25329 8857 25363 8891
rect 5457 8789 5491 8823
rect 12541 8789 12575 8823
rect 17049 8789 17083 8823
rect 23305 8789 23339 8823
rect 24409 8789 24443 8823
rect 5365 8585 5399 8619
rect 9689 8585 9723 8619
rect 11713 8585 11747 8619
rect 14197 8585 14231 8619
rect 25421 8585 25455 8619
rect 6101 8517 6135 8551
rect 9505 8517 9539 8551
rect 9873 8517 9907 8551
rect 12725 8517 12759 8551
rect 17325 8517 17359 8551
rect 23213 8517 23247 8551
rect 23397 8517 23431 8551
rect 23949 8517 23983 8551
rect 5181 8449 5215 8483
rect 5365 8449 5399 8483
rect 5549 8449 5583 8483
rect 6009 8449 6043 8483
rect 6193 8449 6227 8483
rect 6561 8449 6595 8483
rect 8033 8449 8067 8483
rect 9321 8449 9355 8483
rect 9781 8449 9815 8483
rect 9965 8449 9999 8483
rect 11621 8449 11655 8483
rect 12633 8449 12667 8483
rect 12817 8449 12851 8483
rect 14381 8449 14415 8483
rect 14473 8449 14507 8483
rect 14657 8449 14691 8483
rect 14749 8449 14783 8483
rect 17049 8449 17083 8483
rect 17141 8449 17175 8483
rect 18981 8449 19015 8483
rect 19441 8449 19475 8483
rect 19625 8449 19659 8483
rect 19901 8449 19935 8483
rect 20085 8449 20119 8483
rect 20177 8449 20211 8483
rect 22753 8449 22787 8483
rect 23305 8449 23339 8483
rect 23673 8449 23707 8483
rect 6469 8381 6503 8415
rect 7941 8381 7975 8415
rect 8401 8381 8435 8415
rect 19073 8381 19107 8415
rect 6929 8313 6963 8347
rect 19809 8313 19843 8347
rect 23029 8313 23063 8347
rect 23581 8313 23615 8347
rect 5641 8245 5675 8279
rect 16865 8245 16899 8279
rect 17325 8245 17359 8279
rect 19901 8245 19935 8279
rect 20269 8245 20303 8279
rect 22845 8245 22879 8279
rect 5273 8041 5307 8075
rect 6193 8041 6227 8075
rect 10793 8041 10827 8075
rect 13185 8041 13219 8075
rect 13553 8041 13587 8075
rect 15945 8041 15979 8075
rect 16773 8041 16807 8075
rect 17233 8041 17267 8075
rect 19625 8041 19659 8075
rect 20085 8041 20119 8075
rect 21189 8041 21223 8075
rect 22201 8041 22235 8075
rect 23765 8041 23799 8075
rect 24869 8041 24903 8075
rect 15853 7973 15887 8007
rect 21557 7973 21591 8007
rect 24409 7973 24443 8007
rect 4721 7905 4755 7939
rect 5181 7905 5215 7939
rect 5549 7905 5583 7939
rect 5641 7905 5675 7939
rect 16865 7905 16899 7939
rect 19717 7905 19751 7939
rect 20821 7905 20855 7939
rect 23305 7905 23339 7939
rect 4353 7837 4387 7871
rect 4537 7837 4571 7871
rect 4813 7837 4847 7871
rect 5457 7837 5491 7871
rect 5733 7837 5767 7871
rect 6285 7837 6319 7871
rect 9413 7837 9447 7871
rect 9597 7837 9631 7871
rect 12541 7837 12575 7871
rect 12633 7837 12667 7871
rect 12725 7837 12759 7871
rect 12909 7837 12943 7871
rect 13001 7837 13035 7871
rect 15761 7837 15795 7871
rect 15991 7837 16025 7871
rect 16129 7837 16163 7871
rect 17049 7837 17083 7871
rect 17509 7837 17543 7871
rect 17601 7837 17635 7871
rect 17785 7837 17819 7871
rect 17877 7837 17911 7871
rect 18153 7837 18187 7871
rect 18337 7837 18371 7871
rect 18429 7837 18463 7871
rect 18521 7837 18555 7871
rect 18613 7837 18647 7871
rect 18797 7837 18831 7871
rect 18889 7837 18923 7871
rect 19533 7837 19567 7871
rect 19809 7837 19843 7871
rect 19993 7837 20027 7871
rect 20269 7837 20303 7871
rect 20361 7837 20395 7871
rect 20545 7837 20579 7871
rect 20637 7837 20671 7871
rect 20913 7837 20947 7871
rect 22017 7837 22051 7871
rect 22937 7837 22971 7871
rect 23121 7837 23155 7871
rect 23397 7837 23431 7871
rect 24041 7837 24075 7871
rect 24133 7837 24167 7871
rect 25053 7837 25087 7871
rect 4445 7769 4479 7803
rect 12265 7769 12299 7803
rect 13737 7769 13771 7803
rect 16773 7769 16807 7803
rect 21833 7769 21867 7803
rect 24593 7769 24627 7803
rect 9505 7701 9539 7735
rect 13369 7701 13403 7735
rect 13537 7701 13571 7735
rect 17325 7701 17359 7735
rect 17969 7701 18003 7735
rect 19073 7701 19107 7735
rect 19257 7701 19291 7735
rect 22753 7701 22787 7735
rect 23857 7701 23891 7735
rect 4721 7497 4755 7531
rect 7941 7497 7975 7531
rect 8309 7497 8343 7531
rect 8861 7497 8895 7531
rect 12173 7497 12207 7531
rect 12725 7497 12759 7531
rect 14105 7497 14139 7531
rect 14565 7497 14599 7531
rect 14933 7497 14967 7531
rect 17877 7497 17911 7531
rect 18061 7497 18095 7531
rect 18337 7497 18371 7531
rect 20637 7497 20671 7531
rect 22569 7497 22603 7531
rect 23305 7497 23339 7531
rect 25237 7497 25271 7531
rect 9413 7429 9447 7463
rect 10425 7429 10459 7463
rect 10609 7429 10643 7463
rect 10793 7429 10827 7463
rect 11529 7429 11563 7463
rect 15209 7429 15243 7463
rect 15669 7429 15703 7463
rect 20269 7429 20303 7463
rect 23765 7429 23799 7463
rect 4629 7361 4663 7395
rect 4813 7361 4847 7395
rect 5273 7361 5307 7395
rect 5733 7361 5767 7395
rect 6377 7361 6411 7395
rect 6561 7361 6595 7395
rect 8125 7361 8159 7395
rect 8401 7361 8435 7395
rect 8493 7361 8527 7395
rect 8677 7361 8711 7395
rect 9137 7361 9171 7395
rect 9229 7361 9263 7395
rect 9505 7361 9539 7395
rect 9689 7361 9723 7395
rect 9873 7361 9907 7395
rect 9965 7361 9999 7395
rect 10149 7361 10183 7395
rect 10333 7361 10367 7395
rect 11621 7361 11655 7395
rect 11897 7361 11931 7395
rect 13001 7361 13035 7395
rect 13185 7361 13219 7395
rect 13461 7361 13495 7395
rect 13553 7361 13587 7395
rect 13829 7361 13863 7395
rect 13921 7361 13955 7395
rect 14473 7361 14507 7395
rect 14841 7361 14875 7395
rect 15117 7361 15151 7395
rect 15301 7361 15335 7395
rect 15485 7361 15519 7395
rect 15577 7361 15611 7395
rect 15853 7361 15887 7395
rect 15945 7361 15979 7395
rect 16129 7361 16163 7395
rect 16221 7361 16255 7395
rect 16313 7361 16347 7395
rect 16773 7361 16807 7395
rect 16865 7361 16899 7395
rect 17141 7361 17175 7395
rect 17601 7361 17635 7395
rect 17693 7361 17727 7395
rect 18153 7361 18187 7395
rect 18245 7361 18279 7395
rect 19073 7361 19107 7395
rect 19533 7361 19567 7395
rect 20177 7361 20211 7395
rect 20453 7361 20487 7395
rect 20729 7361 20763 7395
rect 20821 7361 20855 7395
rect 21005 7361 21039 7395
rect 21097 7361 21131 7395
rect 21373 7361 21407 7395
rect 21557 7361 21591 7395
rect 21649 7361 21683 7395
rect 21833 7361 21867 7395
rect 22017 7361 22051 7395
rect 22201 7361 22235 7395
rect 22293 7361 22327 7395
rect 22477 7361 22511 7395
rect 23397 7361 23431 7395
rect 23489 7361 23523 7395
rect 5365 7293 5399 7327
rect 5641 7293 5675 7327
rect 6469 7293 6503 7327
rect 11989 7293 12023 7327
rect 13645 7293 13679 7327
rect 14657 7293 14691 7327
rect 16405 7293 16439 7327
rect 16957 7293 16991 7327
rect 17233 7293 17267 7327
rect 17325 7293 17359 7327
rect 19257 7293 19291 7327
rect 19717 7293 19751 7327
rect 6101 7225 6135 7259
rect 17141 7225 17175 7259
rect 21281 7225 21315 7259
rect 22109 7225 22143 7259
rect 4905 7157 4939 7191
rect 13093 7157 13127 7191
rect 13277 7157 13311 7191
rect 14841 7157 14875 7191
rect 21373 7157 21407 7191
rect 8033 6953 8067 6987
rect 9413 6953 9447 6987
rect 9689 6953 9723 6987
rect 12449 6953 12483 6987
rect 13645 6953 13679 6987
rect 15025 6953 15059 6987
rect 15209 6953 15243 6987
rect 15301 6953 15335 6987
rect 15945 6953 15979 6987
rect 20342 6953 20376 6987
rect 21833 6953 21867 6987
rect 8125 6885 8159 6919
rect 11897 6885 11931 6919
rect 5549 6817 5583 6851
rect 7665 6817 7699 6851
rect 9045 6817 9079 6851
rect 14197 6817 14231 6851
rect 17601 6817 17635 6851
rect 19073 6817 19107 6851
rect 20085 6817 20119 6851
rect 5641 6749 5675 6783
rect 7573 6749 7607 6783
rect 8585 6749 8619 6783
rect 8769 6749 8803 6783
rect 9137 6749 9171 6783
rect 9597 6749 9631 6783
rect 9781 6749 9815 6783
rect 10149 6749 10183 6783
rect 10333 6749 10367 6783
rect 12081 6749 12115 6783
rect 12173 6749 12207 6783
rect 12633 6749 12667 6783
rect 12725 6749 12759 6783
rect 12909 6749 12943 6783
rect 13001 6749 13035 6783
rect 13277 6749 13311 6783
rect 13553 6749 13587 6783
rect 13645 6749 13679 6783
rect 13921 6749 13955 6783
rect 14289 6749 14323 6783
rect 14841 6749 14875 6783
rect 14933 6749 14967 6783
rect 15485 6749 15519 6783
rect 15745 6749 15779 6783
rect 15853 6749 15887 6783
rect 17325 6749 17359 6783
rect 23673 6749 23707 6783
rect 24041 6749 24075 6783
rect 8493 6681 8527 6715
rect 11897 6681 11931 6715
rect 13461 6681 13495 6715
rect 13829 6681 13863 6715
rect 15669 6681 15703 6715
rect 6009 6613 6043 6647
rect 7941 6613 7975 6647
rect 8677 6613 8711 6647
rect 10241 6613 10275 6647
rect 13093 6613 13127 6647
rect 14657 6613 14691 6647
rect 18613 6409 18647 6443
rect 27629 6409 27663 6443
rect 11805 6341 11839 6375
rect 16037 6341 16071 6375
rect 17141 6341 17175 6375
rect 8033 6273 8067 6307
rect 8953 6273 8987 6307
rect 11529 6273 11563 6307
rect 13461 6273 13495 6307
rect 13553 6273 13587 6307
rect 16313 6273 16347 6307
rect 16865 6273 16899 6307
rect 27813 6273 27847 6307
rect 8125 6205 8159 6239
rect 8401 6205 8435 6239
rect 8861 6205 8895 6239
rect 9321 6205 9355 6239
rect 13277 6205 13311 6239
rect 14565 6205 14599 6239
rect 8677 5865 8711 5899
rect 27629 5865 27663 5899
rect 8401 5661 8435 5695
rect 8493 5661 8527 5695
rect 8677 5661 8711 5695
rect 27813 5661 27847 5695
rect 6101 2601 6135 2635
rect 9321 2601 9355 2635
rect 5917 2397 5951 2431
rect 9137 2397 9171 2431
<< metal1 >>
rect 1104 28858 28152 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 28152 28858
rect 1104 28784 28152 28806
rect 11790 28704 11796 28756
rect 11848 28704 11854 28756
rect 12342 28704 12348 28756
rect 12400 28744 12406 28756
rect 12437 28747 12495 28753
rect 12437 28744 12449 28747
rect 12400 28716 12449 28744
rect 12400 28704 12406 28716
rect 12437 28713 12449 28716
rect 12483 28713 12495 28747
rect 12437 28707 12495 28713
rect 13078 28704 13084 28756
rect 13136 28704 13142 28756
rect 13722 28704 13728 28756
rect 13780 28704 13786 28756
rect 14366 28704 14372 28756
rect 14424 28704 14430 28756
rect 15010 28704 15016 28756
rect 15068 28704 15074 28756
rect 15654 28704 15660 28756
rect 15712 28704 15718 28756
rect 16298 28704 16304 28756
rect 16356 28704 16362 28756
rect 16942 28704 16948 28756
rect 17000 28704 17006 28756
rect 17586 28704 17592 28756
rect 17644 28704 17650 28756
rect 18230 28704 18236 28756
rect 18288 28704 18294 28756
rect 18874 28704 18880 28756
rect 18932 28704 18938 28756
rect 19610 28704 19616 28756
rect 19668 28704 19674 28756
rect 20254 28704 20260 28756
rect 20312 28704 20318 28756
rect 20530 28704 20536 28756
rect 20588 28744 20594 28756
rect 20901 28747 20959 28753
rect 20901 28744 20913 28747
rect 20588 28716 20913 28744
rect 20588 28704 20594 28716
rect 20901 28713 20913 28716
rect 20947 28713 20959 28747
rect 20901 28707 20959 28713
rect 21542 28704 21548 28756
rect 21600 28704 21606 28756
rect 22002 28704 22008 28756
rect 22060 28744 22066 28756
rect 22097 28747 22155 28753
rect 22097 28744 22109 28747
rect 22060 28716 22109 28744
rect 22060 28704 22066 28716
rect 22097 28713 22109 28716
rect 22143 28713 22155 28747
rect 22097 28707 22155 28713
rect 22830 28704 22836 28756
rect 22888 28704 22894 28756
rect 23382 28704 23388 28756
rect 23440 28744 23446 28756
rect 23477 28747 23535 28753
rect 23477 28744 23489 28747
rect 23440 28716 23489 28744
rect 23440 28704 23446 28716
rect 23477 28713 23489 28716
rect 23523 28713 23535 28747
rect 23477 28707 23535 28713
rect 24118 28704 24124 28756
rect 24176 28704 24182 28756
rect 24762 28704 24768 28756
rect 24820 28704 24826 28756
rect 25406 28704 25412 28756
rect 25464 28704 25470 28756
rect 26050 28704 26056 28756
rect 26108 28704 26114 28756
rect 26694 28704 26700 28756
rect 26752 28704 26758 28756
rect 27338 28704 27344 28756
rect 27396 28704 27402 28756
rect 27709 28747 27767 28753
rect 27709 28713 27721 28747
rect 27755 28744 27767 28747
rect 27798 28744 27804 28756
rect 27755 28716 27804 28744
rect 27755 28713 27767 28716
rect 27709 28707 27767 28713
rect 27798 28704 27804 28716
rect 27856 28704 27862 28756
rect 18138 28676 18144 28688
rect 14568 28648 18144 28676
rect 11974 28500 11980 28552
rect 12032 28500 12038 28552
rect 12621 28543 12679 28549
rect 12621 28509 12633 28543
rect 12667 28509 12679 28543
rect 12621 28503 12679 28509
rect 12636 28404 12664 28503
rect 13262 28500 13268 28552
rect 13320 28500 13326 28552
rect 14568 28549 14596 28648
rect 18138 28636 18144 28648
rect 18196 28636 18202 28688
rect 17954 28608 17960 28620
rect 15120 28580 17960 28608
rect 13909 28543 13967 28549
rect 13909 28509 13921 28543
rect 13955 28509 13967 28543
rect 13909 28503 13967 28509
rect 14553 28543 14611 28549
rect 14553 28509 14565 28543
rect 14599 28509 14611 28543
rect 14553 28503 14611 28509
rect 13924 28472 13952 28503
rect 15120 28472 15148 28580
rect 17954 28568 17960 28580
rect 18012 28568 18018 28620
rect 19978 28608 19984 28620
rect 18340 28580 19984 28608
rect 15197 28543 15255 28549
rect 15197 28509 15209 28543
rect 15243 28509 15255 28543
rect 15197 28503 15255 28509
rect 13924 28444 15148 28472
rect 15212 28472 15240 28503
rect 15838 28500 15844 28552
rect 15896 28500 15902 28552
rect 16485 28543 16543 28549
rect 16485 28509 16497 28543
rect 16531 28540 16543 28543
rect 16942 28540 16948 28552
rect 16531 28512 16948 28540
rect 16531 28509 16543 28512
rect 16485 28503 16543 28509
rect 16942 28500 16948 28512
rect 17000 28500 17006 28552
rect 17126 28500 17132 28552
rect 17184 28500 17190 28552
rect 17773 28543 17831 28549
rect 17773 28509 17785 28543
rect 17819 28540 17831 28543
rect 17862 28540 17868 28552
rect 17819 28512 17868 28540
rect 17819 28509 17831 28512
rect 17773 28503 17831 28509
rect 17862 28500 17868 28512
rect 17920 28500 17926 28552
rect 17402 28472 17408 28484
rect 15212 28444 17408 28472
rect 17402 28432 17408 28444
rect 17460 28432 17466 28484
rect 18340 28472 18368 28580
rect 19978 28568 19984 28580
rect 20036 28568 20042 28620
rect 18417 28543 18475 28549
rect 18417 28509 18429 28543
rect 18463 28509 18475 28543
rect 18417 28503 18475 28509
rect 17788 28444 18368 28472
rect 18432 28472 18460 28503
rect 19058 28500 19064 28552
rect 19116 28500 19122 28552
rect 19426 28500 19432 28552
rect 19484 28500 19490 28552
rect 19886 28500 19892 28552
rect 19944 28540 19950 28552
rect 20073 28543 20131 28549
rect 20073 28540 20085 28543
rect 19944 28512 20085 28540
rect 19944 28500 19950 28512
rect 20073 28509 20085 28512
rect 20119 28509 20131 28543
rect 20073 28503 20131 28509
rect 20438 28500 20444 28552
rect 20496 28540 20502 28552
rect 20717 28543 20775 28549
rect 20717 28540 20729 28543
rect 20496 28512 20729 28540
rect 20496 28500 20502 28512
rect 20717 28509 20729 28512
rect 20763 28509 20775 28543
rect 20717 28503 20775 28509
rect 21358 28500 21364 28552
rect 21416 28500 21422 28552
rect 22278 28500 22284 28552
rect 22336 28500 22342 28552
rect 22646 28500 22652 28552
rect 22704 28500 22710 28552
rect 23290 28500 23296 28552
rect 23348 28500 23354 28552
rect 23934 28500 23940 28552
rect 23992 28500 23998 28552
rect 24578 28500 24584 28552
rect 24636 28500 24642 28552
rect 24946 28500 24952 28552
rect 25004 28540 25010 28552
rect 25225 28543 25283 28549
rect 25225 28540 25237 28543
rect 25004 28512 25237 28540
rect 25004 28500 25010 28512
rect 25225 28509 25237 28512
rect 25271 28509 25283 28543
rect 25225 28503 25283 28509
rect 25866 28500 25872 28552
rect 25924 28500 25930 28552
rect 26050 28500 26056 28552
rect 26108 28540 26114 28552
rect 26513 28543 26571 28549
rect 26513 28540 26525 28543
rect 26108 28512 26525 28540
rect 26108 28500 26114 28512
rect 26513 28509 26525 28512
rect 26559 28509 26571 28543
rect 26513 28503 26571 28509
rect 26786 28500 26792 28552
rect 26844 28540 26850 28552
rect 27157 28543 27215 28549
rect 27157 28540 27169 28543
rect 26844 28512 27169 28540
rect 26844 28500 26850 28512
rect 27157 28509 27169 28512
rect 27203 28509 27215 28543
rect 27157 28503 27215 28509
rect 27525 28543 27583 28549
rect 27525 28509 27537 28543
rect 27571 28509 27583 28543
rect 27525 28503 27583 28509
rect 21450 28472 21456 28484
rect 18432 28444 21456 28472
rect 17788 28416 17816 28444
rect 21450 28432 21456 28444
rect 21508 28432 21514 28484
rect 26142 28432 26148 28484
rect 26200 28472 26206 28484
rect 27540 28472 27568 28503
rect 26200 28444 27568 28472
rect 26200 28432 26206 28444
rect 17218 28404 17224 28416
rect 12636 28376 17224 28404
rect 17218 28364 17224 28376
rect 17276 28364 17282 28416
rect 17770 28364 17776 28416
rect 17828 28364 17834 28416
rect 18690 28364 18696 28416
rect 18748 28404 18754 28416
rect 20070 28404 20076 28416
rect 18748 28376 20076 28404
rect 18748 28364 18754 28376
rect 20070 28364 20076 28376
rect 20128 28364 20134 28416
rect 1104 28314 28152 28336
rect 1104 28262 4874 28314
rect 4926 28262 4938 28314
rect 4990 28262 5002 28314
rect 5054 28262 5066 28314
rect 5118 28262 5130 28314
rect 5182 28262 28152 28314
rect 1104 28240 28152 28262
rect 17126 28160 17132 28212
rect 17184 28200 17190 28212
rect 18969 28203 19027 28209
rect 18969 28200 18981 28203
rect 17184 28172 18981 28200
rect 17184 28160 17190 28172
rect 18969 28169 18981 28172
rect 19015 28169 19027 28203
rect 18969 28163 19027 28169
rect 19058 28160 19064 28212
rect 19116 28200 19122 28212
rect 20165 28203 20223 28209
rect 20165 28200 20177 28203
rect 19116 28172 20177 28200
rect 19116 28160 19122 28172
rect 20165 28169 20177 28172
rect 20211 28169 20223 28203
rect 20165 28163 20223 28169
rect 20438 28160 20444 28212
rect 20496 28160 20502 28212
rect 24946 28160 24952 28212
rect 25004 28160 25010 28212
rect 27709 28203 27767 28209
rect 27709 28169 27721 28203
rect 27755 28200 27767 28203
rect 28718 28200 28724 28212
rect 27755 28172 28724 28200
rect 27755 28169 27767 28172
rect 27709 28163 27767 28169
rect 28718 28160 28724 28172
rect 28776 28160 28782 28212
rect 10336 28104 11284 28132
rect 7466 27956 7472 28008
rect 7524 27996 7530 28008
rect 10336 28005 10364 28104
rect 11054 28024 11060 28076
rect 11112 28073 11118 28076
rect 11256 28073 11284 28104
rect 13262 28092 13268 28144
rect 13320 28132 13326 28144
rect 19613 28135 19671 28141
rect 19613 28132 19625 28135
rect 13320 28104 19625 28132
rect 13320 28092 13326 28104
rect 19613 28101 19625 28104
rect 19659 28101 19671 28135
rect 19613 28095 19671 28101
rect 20180 28104 20576 28132
rect 11112 28067 11145 28073
rect 11133 28033 11145 28067
rect 11112 28027 11145 28033
rect 11241 28067 11299 28073
rect 11241 28033 11253 28067
rect 11287 28064 11299 28067
rect 11698 28064 11704 28076
rect 11287 28036 11704 28064
rect 11287 28033 11299 28036
rect 11241 28027 11299 28033
rect 11112 28024 11118 28027
rect 11698 28024 11704 28036
rect 11756 28024 11762 28076
rect 11974 28024 11980 28076
rect 12032 28064 12038 28076
rect 18598 28064 18604 28076
rect 12032 28036 18604 28064
rect 12032 28024 12038 28036
rect 18598 28024 18604 28036
rect 18656 28024 18662 28076
rect 18690 28024 18696 28076
rect 18748 28024 18754 28076
rect 19153 28067 19211 28073
rect 19153 28033 19165 28067
rect 19199 28033 19211 28067
rect 19153 28027 19211 28033
rect 19245 28067 19303 28073
rect 19245 28033 19257 28067
rect 19291 28033 19303 28067
rect 19245 28027 19303 28033
rect 19337 28067 19395 28073
rect 19337 28033 19349 28067
rect 19383 28064 19395 28067
rect 19518 28064 19524 28076
rect 19383 28036 19524 28064
rect 19383 28033 19395 28036
rect 19337 28027 19395 28033
rect 10321 27999 10379 28005
rect 10321 27996 10333 27999
rect 7524 27968 10333 27996
rect 7524 27956 7530 27968
rect 10321 27965 10333 27968
rect 10367 27965 10379 27999
rect 10321 27959 10379 27965
rect 15838 27956 15844 28008
rect 15896 27996 15902 28008
rect 19058 27996 19064 28008
rect 15896 27968 19064 27996
rect 15896 27956 15902 27968
rect 19058 27956 19064 27968
rect 19116 27956 19122 28008
rect 19168 27940 19196 28027
rect 19260 27996 19288 28027
rect 19518 28024 19524 28036
rect 19576 28024 19582 28076
rect 19797 28067 19855 28073
rect 19797 28033 19809 28067
rect 19843 28033 19855 28067
rect 19797 28027 19855 28033
rect 19610 27996 19616 28008
rect 19260 27968 19616 27996
rect 19610 27956 19616 27968
rect 19668 27956 19674 28008
rect 10686 27888 10692 27940
rect 10744 27888 10750 27940
rect 10781 27931 10839 27937
rect 10781 27897 10793 27931
rect 10827 27928 10839 27931
rect 11146 27928 11152 27940
rect 10827 27900 11152 27928
rect 10827 27897 10839 27900
rect 10781 27891 10839 27897
rect 11146 27888 11152 27900
rect 11204 27888 11210 27940
rect 18046 27888 18052 27940
rect 18104 27928 18110 27940
rect 19150 27928 19156 27940
rect 18104 27900 19156 27928
rect 18104 27888 18110 27900
rect 19150 27888 19156 27900
rect 19208 27888 19214 27940
rect 19521 27931 19579 27937
rect 19521 27897 19533 27931
rect 19567 27928 19579 27931
rect 19702 27928 19708 27940
rect 19567 27900 19708 27928
rect 19567 27897 19579 27900
rect 19521 27891 19579 27897
rect 19702 27888 19708 27900
rect 19760 27888 19766 27940
rect 19812 27928 19840 28027
rect 20070 28024 20076 28076
rect 20128 28073 20134 28076
rect 20128 28064 20137 28073
rect 20180 28064 20208 28104
rect 20128 28036 20208 28064
rect 20257 28067 20315 28073
rect 20128 28027 20137 28036
rect 20257 28033 20269 28067
rect 20303 28033 20315 28067
rect 20257 28027 20315 28033
rect 20128 28024 20134 28027
rect 19978 27956 19984 28008
rect 20036 27956 20042 28008
rect 20272 27996 20300 28027
rect 20346 28024 20352 28076
rect 20404 28024 20410 28076
rect 20548 28073 20576 28104
rect 21652 28104 24900 28132
rect 21652 28076 21680 28104
rect 20533 28067 20591 28073
rect 20533 28033 20545 28067
rect 20579 28064 20591 28067
rect 20579 28036 21588 28064
rect 20579 28033 20591 28036
rect 20533 28027 20591 28033
rect 21082 27996 21088 28008
rect 20272 27968 21088 27996
rect 21082 27956 21088 27968
rect 21140 27956 21146 28008
rect 20990 27928 20996 27940
rect 19812 27900 20996 27928
rect 20990 27888 20996 27900
rect 21048 27888 21054 27940
rect 21560 27928 21588 28036
rect 21634 28024 21640 28076
rect 21692 28024 21698 28076
rect 22005 28067 22063 28073
rect 22005 28033 22017 28067
rect 22051 28033 22063 28067
rect 22005 28027 22063 28033
rect 22020 27996 22048 28027
rect 22094 28024 22100 28076
rect 22152 28064 22158 28076
rect 22189 28067 22247 28073
rect 22189 28064 22201 28067
rect 22152 28036 22201 28064
rect 22152 28024 22158 28036
rect 22189 28033 22201 28036
rect 22235 28064 22247 28067
rect 23382 28064 23388 28076
rect 22235 28036 23388 28064
rect 22235 28033 22247 28036
rect 22189 28027 22247 28033
rect 23382 28024 23388 28036
rect 23440 28024 23446 28076
rect 24872 28073 24900 28104
rect 24857 28067 24915 28073
rect 24857 28033 24869 28067
rect 24903 28064 24915 28067
rect 24946 28064 24952 28076
rect 24903 28036 24952 28064
rect 24903 28033 24915 28036
rect 24857 28027 24915 28033
rect 24946 28024 24952 28036
rect 25004 28024 25010 28076
rect 25038 28024 25044 28076
rect 25096 28024 25102 28076
rect 27154 28024 27160 28076
rect 27212 28024 27218 28076
rect 27525 28067 27583 28073
rect 27525 28033 27537 28067
rect 27571 28033 27583 28067
rect 27525 28027 27583 28033
rect 22370 27996 22376 28008
rect 22020 27968 22376 27996
rect 22370 27956 22376 27968
rect 22428 27956 22434 28008
rect 25406 27956 25412 28008
rect 25464 27996 25470 28008
rect 27540 27996 27568 28027
rect 25464 27968 27568 27996
rect 25464 27956 25470 27968
rect 24026 27928 24032 27940
rect 21560 27900 24032 27928
rect 24026 27888 24032 27900
rect 24084 27928 24090 27940
rect 26234 27928 26240 27940
rect 24084 27900 26240 27928
rect 24084 27888 24090 27900
rect 26234 27888 26240 27900
rect 26292 27888 26298 27940
rect 27341 27931 27399 27937
rect 27341 27897 27353 27931
rect 27387 27928 27399 27931
rect 27982 27928 27988 27940
rect 27387 27900 27988 27928
rect 27387 27897 27399 27900
rect 27341 27891 27399 27897
rect 27982 27888 27988 27900
rect 28040 27888 28046 27940
rect 11057 27863 11115 27869
rect 11057 27829 11069 27863
rect 11103 27860 11115 27863
rect 11238 27860 11244 27872
rect 11103 27832 11244 27860
rect 11103 27829 11115 27832
rect 11057 27823 11115 27829
rect 11238 27820 11244 27832
rect 11296 27820 11302 27872
rect 18601 27863 18659 27869
rect 18601 27829 18613 27863
rect 18647 27860 18659 27863
rect 18782 27860 18788 27872
rect 18647 27832 18788 27860
rect 18647 27829 18659 27832
rect 18601 27823 18659 27829
rect 18782 27820 18788 27832
rect 18840 27820 18846 27872
rect 19168 27860 19196 27888
rect 21542 27860 21548 27872
rect 19168 27832 21548 27860
rect 21542 27820 21548 27832
rect 21600 27820 21606 27872
rect 22094 27820 22100 27872
rect 22152 27860 22158 27872
rect 22189 27863 22247 27869
rect 22189 27860 22201 27863
rect 22152 27832 22201 27860
rect 22152 27820 22158 27832
rect 22189 27829 22201 27832
rect 22235 27829 22247 27863
rect 22189 27823 22247 27829
rect 1104 27770 28152 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 28152 27770
rect 1104 27696 28152 27718
rect 2774 27616 2780 27668
rect 2832 27656 2838 27668
rect 6825 27659 6883 27665
rect 2832 27628 6592 27656
rect 2832 27616 2838 27628
rect 3142 27548 3148 27600
rect 3200 27588 3206 27600
rect 3200 27560 5212 27588
rect 3200 27548 3206 27560
rect 4614 27480 4620 27532
rect 4672 27520 4678 27532
rect 5077 27523 5135 27529
rect 5077 27520 5089 27523
rect 4672 27492 5089 27520
rect 4672 27480 4678 27492
rect 5077 27489 5089 27492
rect 5123 27489 5135 27523
rect 5184 27528 5212 27560
rect 5442 27548 5448 27600
rect 5500 27588 5506 27600
rect 5500 27560 6224 27588
rect 5500 27548 5506 27560
rect 5264 27528 5322 27529
rect 5184 27523 5386 27528
rect 5184 27500 5276 27523
rect 5077 27483 5135 27489
rect 5264 27489 5276 27500
rect 5310 27520 5386 27523
rect 5718 27520 5724 27532
rect 5310 27500 5724 27520
rect 5310 27489 5322 27500
rect 5358 27492 5724 27500
rect 5264 27483 5322 27489
rect 5718 27480 5724 27492
rect 5776 27480 5782 27532
rect 6196 27520 6224 27560
rect 6196 27492 6316 27520
rect 2038 27412 2044 27464
rect 2096 27452 2102 27464
rect 4985 27455 5043 27461
rect 4985 27452 4997 27455
rect 2096 27424 4997 27452
rect 2096 27412 2102 27424
rect 4985 27421 4997 27424
rect 5031 27452 5043 27455
rect 5166 27452 5172 27464
rect 5031 27424 5172 27452
rect 5031 27421 5043 27424
rect 4985 27415 5043 27421
rect 5166 27412 5172 27424
rect 5224 27412 5230 27464
rect 5353 27455 5411 27461
rect 5353 27421 5365 27455
rect 5399 27452 5411 27455
rect 5537 27455 5595 27461
rect 5399 27424 5488 27452
rect 5399 27421 5411 27424
rect 5353 27415 5411 27421
rect 5460 27384 5488 27424
rect 5537 27421 5549 27455
rect 5583 27452 5595 27455
rect 5813 27455 5871 27461
rect 5813 27452 5825 27455
rect 5583 27424 5825 27452
rect 5583 27421 5595 27424
rect 5537 27415 5595 27421
rect 5813 27421 5825 27424
rect 5859 27452 5871 27455
rect 5902 27452 5908 27464
rect 5859 27424 5908 27452
rect 5859 27421 5871 27424
rect 5813 27415 5871 27421
rect 5902 27412 5908 27424
rect 5960 27412 5966 27464
rect 5994 27412 6000 27464
rect 6052 27412 6058 27464
rect 6089 27455 6147 27461
rect 6089 27421 6101 27455
rect 6135 27421 6147 27455
rect 6089 27415 6147 27421
rect 5626 27384 5632 27396
rect 5460 27356 5632 27384
rect 5626 27344 5632 27356
rect 5684 27344 5690 27396
rect 5718 27344 5724 27396
rect 5776 27384 5782 27396
rect 6104 27384 6132 27415
rect 6178 27412 6184 27464
rect 6236 27412 6242 27464
rect 6288 27461 6316 27492
rect 6564 27461 6592 27628
rect 6825 27625 6837 27659
rect 6871 27656 6883 27659
rect 6914 27656 6920 27668
rect 6871 27628 6920 27656
rect 6871 27625 6883 27628
rect 6825 27619 6883 27625
rect 6914 27616 6920 27628
rect 6972 27616 6978 27668
rect 10318 27616 10324 27668
rect 10376 27616 10382 27668
rect 10428 27628 10824 27656
rect 6730 27548 6736 27600
rect 6788 27588 6794 27600
rect 7466 27588 7472 27600
rect 6788 27560 7472 27588
rect 6788 27548 6794 27560
rect 7466 27548 7472 27560
rect 7524 27548 7530 27600
rect 10428 27588 10456 27628
rect 9968 27560 10456 27588
rect 6641 27523 6699 27529
rect 6641 27489 6653 27523
rect 6687 27520 6699 27523
rect 7009 27523 7067 27529
rect 7009 27520 7021 27523
rect 6687 27492 7021 27520
rect 6687 27489 6699 27492
rect 6641 27483 6699 27489
rect 7009 27489 7021 27492
rect 7055 27489 7067 27523
rect 9968 27520 9996 27560
rect 10502 27548 10508 27600
rect 10560 27588 10566 27600
rect 10689 27591 10747 27597
rect 10689 27588 10701 27591
rect 10560 27560 10701 27588
rect 10560 27548 10566 27560
rect 10689 27557 10701 27560
rect 10735 27557 10747 27591
rect 10796 27588 10824 27628
rect 11054 27616 11060 27668
rect 11112 27656 11118 27668
rect 18141 27659 18199 27665
rect 18141 27656 18153 27659
rect 11112 27628 11836 27656
rect 11112 27616 11118 27628
rect 10962 27588 10968 27600
rect 10796 27560 10968 27588
rect 10689 27551 10747 27557
rect 10962 27548 10968 27560
rect 11020 27588 11026 27600
rect 11020 27560 11468 27588
rect 11020 27548 11026 27560
rect 7009 27483 7067 27489
rect 7300 27492 9996 27520
rect 6273 27455 6331 27461
rect 6273 27421 6285 27455
rect 6319 27421 6331 27455
rect 6273 27415 6331 27421
rect 6549 27455 6607 27461
rect 6549 27421 6561 27455
rect 6595 27452 6607 27455
rect 6822 27452 6828 27464
rect 6595 27424 6828 27452
rect 6595 27421 6607 27424
rect 6549 27415 6607 27421
rect 6288 27384 6316 27415
rect 6822 27412 6828 27424
rect 6880 27412 6886 27464
rect 7193 27433 7251 27439
rect 7193 27430 7205 27433
rect 7116 27402 7205 27430
rect 7116 27384 7144 27402
rect 7193 27399 7205 27402
rect 7239 27430 7251 27433
rect 7300 27430 7328 27492
rect 7239 27402 7328 27430
rect 7466 27412 7472 27464
rect 7524 27412 7530 27464
rect 7650 27412 7656 27464
rect 7708 27452 7714 27464
rect 9968 27461 9996 27492
rect 10336 27492 11192 27520
rect 10336 27461 10364 27492
rect 9493 27455 9551 27461
rect 9324 27452 9444 27454
rect 9493 27452 9505 27455
rect 7708 27426 9505 27452
rect 7708 27424 9352 27426
rect 9416 27424 9505 27426
rect 7708 27412 7714 27424
rect 9493 27421 9505 27424
rect 9539 27421 9551 27455
rect 9493 27415 9551 27421
rect 9953 27455 10011 27461
rect 9953 27421 9965 27455
rect 9999 27421 10011 27455
rect 9953 27415 10011 27421
rect 10321 27455 10379 27461
rect 10321 27421 10333 27455
rect 10367 27421 10379 27455
rect 10321 27415 10379 27421
rect 10594 27412 10600 27464
rect 10652 27412 10658 27464
rect 10778 27412 10784 27464
rect 10836 27412 10842 27464
rect 11164 27461 11192 27492
rect 11149 27455 11207 27461
rect 11149 27421 11161 27455
rect 11195 27452 11207 27455
rect 11238 27452 11244 27464
rect 11195 27424 11244 27452
rect 11195 27421 11207 27424
rect 11149 27415 11207 27421
rect 11238 27412 11244 27424
rect 11296 27412 11302 27464
rect 11440 27461 11468 27560
rect 11808 27520 11836 27628
rect 17880 27628 18153 27656
rect 16942 27548 16948 27600
rect 17000 27548 17006 27600
rect 17218 27548 17224 27600
rect 17276 27548 17282 27600
rect 17770 27548 17776 27600
rect 17828 27588 17834 27600
rect 17880 27588 17908 27628
rect 18141 27625 18153 27628
rect 18187 27625 18199 27659
rect 18141 27619 18199 27625
rect 18230 27616 18236 27668
rect 18288 27656 18294 27668
rect 18782 27656 18788 27668
rect 18288 27628 18788 27656
rect 18288 27616 18294 27628
rect 18782 27616 18788 27628
rect 18840 27656 18846 27668
rect 19242 27656 19248 27668
rect 18840 27628 19248 27656
rect 18840 27616 18846 27628
rect 19242 27616 19248 27628
rect 19300 27616 19306 27668
rect 19886 27616 19892 27668
rect 19944 27616 19950 27668
rect 20070 27616 20076 27668
rect 20128 27616 20134 27668
rect 20806 27616 20812 27668
rect 20864 27616 20870 27668
rect 21008 27628 21312 27656
rect 17828 27560 17908 27588
rect 17828 27548 17834 27560
rect 18598 27548 18604 27600
rect 18656 27548 18662 27600
rect 21008 27588 21036 27628
rect 18800 27560 21036 27588
rect 18800 27532 18828 27560
rect 21082 27548 21088 27600
rect 21140 27548 21146 27600
rect 17497 27523 17555 27529
rect 17497 27520 17509 27523
rect 11808 27492 11928 27520
rect 11900 27464 11928 27492
rect 17236 27492 17509 27520
rect 11425 27455 11483 27461
rect 11425 27421 11437 27455
rect 11471 27421 11483 27455
rect 11425 27415 11483 27421
rect 11698 27412 11704 27464
rect 11756 27461 11762 27464
rect 11756 27455 11789 27461
rect 11777 27421 11789 27455
rect 11756 27415 11789 27421
rect 11756 27412 11762 27415
rect 11882 27412 11888 27464
rect 11940 27412 11946 27464
rect 16942 27412 16948 27464
rect 17000 27412 17006 27464
rect 17236 27461 17264 27492
rect 17497 27489 17509 27492
rect 17543 27489 17555 27523
rect 18690 27520 18696 27532
rect 17497 27483 17555 27489
rect 17696 27492 18696 27520
rect 17129 27455 17187 27461
rect 17129 27421 17141 27455
rect 17175 27452 17187 27455
rect 17221 27455 17279 27461
rect 17221 27452 17233 27455
rect 17175 27424 17233 27452
rect 17175 27421 17187 27424
rect 17129 27415 17187 27421
rect 17221 27421 17233 27424
rect 17267 27421 17279 27455
rect 17221 27415 17279 27421
rect 17405 27455 17463 27461
rect 17405 27421 17417 27455
rect 17451 27452 17463 27455
rect 17696 27452 17724 27492
rect 18690 27480 18696 27492
rect 18748 27480 18754 27532
rect 18782 27480 18788 27532
rect 18840 27480 18846 27532
rect 18984 27492 20300 27520
rect 17451 27424 17724 27452
rect 17772 27455 17830 27461
rect 17451 27421 17463 27424
rect 17405 27415 17463 27421
rect 17772 27421 17784 27455
rect 17818 27421 17830 27455
rect 17772 27415 17830 27421
rect 17865 27455 17923 27461
rect 17865 27421 17877 27455
rect 17911 27452 17923 27455
rect 18506 27452 18512 27464
rect 17911 27424 18512 27452
rect 17911 27421 17923 27424
rect 17865 27415 17923 27421
rect 7239 27399 7251 27402
rect 7193 27393 7251 27399
rect 5776 27356 6224 27384
rect 6288 27356 7144 27384
rect 9677 27387 9735 27393
rect 5776 27344 5782 27356
rect 5261 27319 5319 27325
rect 5261 27285 5273 27319
rect 5307 27316 5319 27319
rect 5350 27316 5356 27328
rect 5307 27288 5356 27316
rect 5307 27285 5319 27288
rect 5261 27279 5319 27285
rect 5350 27276 5356 27288
rect 5408 27276 5414 27328
rect 5442 27276 5448 27328
rect 5500 27276 5506 27328
rect 5534 27276 5540 27328
rect 5592 27316 5598 27328
rect 5813 27319 5871 27325
rect 5813 27316 5825 27319
rect 5592 27288 5825 27316
rect 5592 27276 5598 27288
rect 5813 27285 5825 27288
rect 5859 27285 5871 27319
rect 6196 27316 6224 27356
rect 9677 27353 9689 27387
rect 9723 27384 9735 27387
rect 9861 27387 9919 27393
rect 9723 27356 9757 27384
rect 9723 27353 9735 27356
rect 9677 27347 9735 27353
rect 9861 27353 9873 27387
rect 9907 27384 9919 27387
rect 10796 27384 10824 27412
rect 9907 27356 10824 27384
rect 17788 27384 17816 27415
rect 18506 27412 18512 27424
rect 18564 27452 18570 27464
rect 18984 27452 19012 27492
rect 20272 27464 20300 27492
rect 18564 27424 19012 27452
rect 18564 27412 18570 27424
rect 18984 27393 19012 27424
rect 19242 27412 19248 27464
rect 19300 27452 19306 27464
rect 19429 27455 19487 27461
rect 19429 27452 19441 27455
rect 19300 27424 19441 27452
rect 19300 27412 19306 27424
rect 19429 27421 19441 27424
rect 19475 27421 19487 27455
rect 19429 27415 19487 27421
rect 19521 27455 19579 27461
rect 19521 27421 19533 27455
rect 19567 27452 19579 27455
rect 19610 27452 19616 27464
rect 19567 27424 19616 27452
rect 19567 27421 19579 27424
rect 19521 27415 19579 27421
rect 19610 27412 19616 27424
rect 19668 27412 19674 27464
rect 20254 27412 20260 27464
rect 20312 27452 20318 27464
rect 20441 27455 20499 27461
rect 20441 27452 20453 27455
rect 20312 27424 20453 27452
rect 20312 27412 20318 27424
rect 20441 27421 20453 27424
rect 20487 27421 20499 27455
rect 20441 27415 20499 27421
rect 20533 27455 20591 27461
rect 20533 27421 20545 27455
rect 20579 27421 20591 27455
rect 20533 27415 20591 27421
rect 18969 27387 19027 27393
rect 17788 27356 18368 27384
rect 9907 27353 9919 27356
rect 9861 27347 9919 27353
rect 6730 27316 6736 27328
rect 6196 27288 6736 27316
rect 5813 27279 5871 27285
rect 6730 27276 6736 27288
rect 6788 27276 6794 27328
rect 6822 27276 6828 27328
rect 6880 27316 6886 27328
rect 9692 27316 9720 27347
rect 18340 27328 18368 27356
rect 18969 27353 18981 27387
rect 19015 27353 19027 27387
rect 18969 27347 19027 27353
rect 19150 27344 19156 27396
rect 19208 27384 19214 27396
rect 19208 27356 19748 27384
rect 19208 27344 19214 27356
rect 10318 27316 10324 27328
rect 6880 27288 10324 27316
rect 6880 27276 6886 27288
rect 10318 27276 10324 27288
rect 10376 27276 10382 27328
rect 10410 27276 10416 27328
rect 10468 27316 10474 27328
rect 10505 27319 10563 27325
rect 10505 27316 10517 27319
rect 10468 27288 10517 27316
rect 10468 27276 10474 27288
rect 10505 27285 10517 27288
rect 10551 27285 10563 27319
rect 10505 27279 10563 27285
rect 10594 27276 10600 27328
rect 10652 27316 10658 27328
rect 11517 27319 11575 27325
rect 11517 27316 11529 27319
rect 10652 27288 11529 27316
rect 10652 27276 10658 27288
rect 11517 27285 11529 27288
rect 11563 27316 11575 27319
rect 11974 27316 11980 27328
rect 11563 27288 11980 27316
rect 11563 27285 11575 27288
rect 11517 27279 11575 27285
rect 11974 27276 11980 27288
rect 12032 27276 12038 27328
rect 17954 27276 17960 27328
rect 18012 27276 18018 27328
rect 18141 27319 18199 27325
rect 18141 27285 18153 27319
rect 18187 27316 18199 27319
rect 18230 27316 18236 27328
rect 18187 27288 18236 27316
rect 18187 27285 18199 27288
rect 18141 27279 18199 27285
rect 18230 27276 18236 27288
rect 18288 27276 18294 27328
rect 18322 27276 18328 27328
rect 18380 27316 18386 27328
rect 18759 27319 18817 27325
rect 18759 27316 18771 27319
rect 18380 27288 18771 27316
rect 18380 27276 18386 27288
rect 18759 27285 18771 27288
rect 18805 27285 18817 27319
rect 18759 27279 18817 27285
rect 19058 27276 19064 27328
rect 19116 27316 19122 27328
rect 19245 27319 19303 27325
rect 19245 27316 19257 27319
rect 19116 27288 19257 27316
rect 19116 27276 19122 27288
rect 19245 27285 19257 27288
rect 19291 27285 19303 27319
rect 19245 27279 19303 27285
rect 19518 27276 19524 27328
rect 19576 27316 19582 27328
rect 19613 27319 19671 27325
rect 19613 27316 19625 27319
rect 19576 27288 19625 27316
rect 19576 27276 19582 27288
rect 19613 27285 19625 27288
rect 19659 27285 19671 27319
rect 19720 27316 19748 27356
rect 19794 27344 19800 27396
rect 19852 27344 19858 27396
rect 20162 27344 20168 27396
rect 20220 27384 20226 27396
rect 20548 27384 20576 27415
rect 20898 27412 20904 27464
rect 20956 27412 20962 27464
rect 21100 27452 21128 27548
rect 21284 27520 21312 27628
rect 21358 27616 21364 27668
rect 21416 27616 21422 27668
rect 22278 27616 22284 27668
rect 22336 27656 22342 27668
rect 22373 27659 22431 27665
rect 22373 27656 22385 27659
rect 22336 27628 22385 27656
rect 22336 27616 22342 27628
rect 22373 27625 22385 27628
rect 22419 27625 22431 27659
rect 22373 27619 22431 27625
rect 23753 27659 23811 27665
rect 23753 27625 23765 27659
rect 23799 27656 23811 27659
rect 23934 27656 23940 27668
rect 23799 27628 23940 27656
rect 23799 27625 23811 27628
rect 23753 27619 23811 27625
rect 23934 27616 23940 27628
rect 23992 27616 23998 27668
rect 24213 27659 24271 27665
rect 24213 27625 24225 27659
rect 24259 27656 24271 27659
rect 24578 27656 24584 27668
rect 24259 27628 24584 27656
rect 24259 27625 24271 27628
rect 24213 27619 24271 27625
rect 24578 27616 24584 27628
rect 24636 27616 24642 27668
rect 24670 27616 24676 27668
rect 24728 27656 24734 27668
rect 24857 27659 24915 27665
rect 24857 27656 24869 27659
rect 24728 27628 24869 27656
rect 24728 27616 24734 27628
rect 24857 27625 24869 27628
rect 24903 27625 24915 27659
rect 24857 27619 24915 27625
rect 25038 27616 25044 27668
rect 25096 27656 25102 27668
rect 25133 27659 25191 27665
rect 25133 27656 25145 27659
rect 25096 27628 25145 27656
rect 25096 27616 25102 27628
rect 25133 27625 25145 27628
rect 25179 27625 25191 27659
rect 25133 27619 25191 27625
rect 25685 27659 25743 27665
rect 25685 27625 25697 27659
rect 25731 27625 25743 27659
rect 25685 27619 25743 27625
rect 21450 27548 21456 27600
rect 21508 27548 21514 27600
rect 22189 27591 22247 27597
rect 22189 27557 22201 27591
rect 22235 27588 22247 27591
rect 22554 27588 22560 27600
rect 22235 27560 22560 27588
rect 22235 27557 22247 27560
rect 22189 27551 22247 27557
rect 22554 27548 22560 27560
rect 22612 27548 22618 27600
rect 25700 27588 25728 27619
rect 25958 27616 25964 27668
rect 26016 27656 26022 27668
rect 26145 27659 26203 27665
rect 26145 27656 26157 27659
rect 26016 27628 26157 27656
rect 26016 27616 26022 27628
rect 26145 27625 26157 27628
rect 26191 27625 26203 27659
rect 26145 27619 26203 27625
rect 26786 27616 26792 27668
rect 26844 27616 26850 27668
rect 27154 27616 27160 27668
rect 27212 27656 27218 27668
rect 27249 27659 27307 27665
rect 27249 27656 27261 27659
rect 27212 27628 27261 27656
rect 27212 27616 27218 27628
rect 27249 27625 27261 27628
rect 27295 27625 27307 27659
rect 27249 27619 27307 27625
rect 24872 27560 25728 27588
rect 24872 27532 24900 27560
rect 21634 27520 21640 27532
rect 21284 27492 21640 27520
rect 21177 27455 21235 27461
rect 21177 27452 21189 27455
rect 21100 27424 21189 27452
rect 21177 27421 21189 27424
rect 21223 27421 21235 27455
rect 21284 27452 21312 27492
rect 21634 27480 21640 27492
rect 21692 27480 21698 27532
rect 21729 27523 21787 27529
rect 21729 27489 21741 27523
rect 21775 27520 21787 27523
rect 22094 27520 22100 27532
rect 21775 27492 22100 27520
rect 21775 27489 21787 27492
rect 21729 27483 21787 27489
rect 22094 27480 22100 27492
rect 22152 27520 22158 27532
rect 22741 27523 22799 27529
rect 22741 27520 22753 27523
rect 22152 27492 22753 27520
rect 22152 27480 22158 27492
rect 22741 27489 22753 27492
rect 22787 27489 22799 27523
rect 22741 27483 22799 27489
rect 24489 27523 24547 27529
rect 24489 27489 24501 27523
rect 24535 27520 24547 27523
rect 24854 27520 24860 27532
rect 24535 27492 24860 27520
rect 24535 27489 24547 27492
rect 24489 27483 24547 27489
rect 24854 27480 24860 27492
rect 24912 27480 24918 27532
rect 25314 27529 25320 27532
rect 25299 27523 25320 27529
rect 25299 27489 25311 27523
rect 25299 27483 25320 27489
rect 25314 27480 25320 27483
rect 25372 27480 25378 27532
rect 25700 27520 25728 27560
rect 25774 27548 25780 27600
rect 25832 27588 25838 27600
rect 25832 27560 26556 27588
rect 25832 27548 25838 27560
rect 25700 27492 26096 27520
rect 21361 27455 21419 27461
rect 21361 27452 21373 27455
rect 21284 27424 21373 27452
rect 21177 27415 21235 27421
rect 21361 27421 21373 27424
rect 21407 27421 21419 27455
rect 21361 27415 21419 27421
rect 21652 27424 22692 27452
rect 20220 27356 20576 27384
rect 20220 27344 20226 27356
rect 20990 27344 20996 27396
rect 21048 27384 21054 27396
rect 21652 27393 21680 27424
rect 21637 27387 21695 27393
rect 21637 27384 21649 27387
rect 21048 27356 21649 27384
rect 21048 27344 21054 27356
rect 21637 27353 21649 27356
rect 21683 27353 21695 27387
rect 21637 27347 21695 27353
rect 22186 27344 22192 27396
rect 22244 27344 22250 27396
rect 22554 27393 22560 27396
rect 22532 27387 22560 27393
rect 22532 27353 22544 27387
rect 22532 27347 22560 27353
rect 22547 27344 22560 27347
rect 22612 27344 22618 27396
rect 22664 27393 22692 27424
rect 23014 27412 23020 27464
rect 23072 27412 23078 27464
rect 23106 27412 23112 27464
rect 23164 27412 23170 27464
rect 23382 27412 23388 27464
rect 23440 27412 23446 27464
rect 24026 27412 24032 27464
rect 24084 27412 24090 27464
rect 24210 27412 24216 27464
rect 24268 27412 24274 27464
rect 24394 27412 24400 27464
rect 24452 27452 24458 27464
rect 24581 27455 24639 27461
rect 24581 27452 24593 27455
rect 24452 27424 24593 27452
rect 24452 27412 24458 27424
rect 24581 27421 24593 27424
rect 24627 27421 24639 27455
rect 24581 27415 24639 27421
rect 22649 27387 22707 27393
rect 22649 27353 22661 27387
rect 22695 27384 22707 27387
rect 23477 27387 23535 27393
rect 23477 27384 23489 27387
rect 22695 27356 23489 27384
rect 22695 27353 22707 27356
rect 22649 27347 22707 27353
rect 23477 27353 23489 27356
rect 23523 27353 23535 27387
rect 23477 27347 23535 27353
rect 23594 27387 23652 27393
rect 23594 27353 23606 27387
rect 23640 27384 23652 27387
rect 23750 27384 23756 27396
rect 23640 27356 23756 27384
rect 23640 27353 23652 27356
rect 23594 27347 23652 27353
rect 20073 27319 20131 27325
rect 20073 27316 20085 27319
rect 19720 27288 20085 27316
rect 19613 27279 19671 27285
rect 20073 27285 20085 27288
rect 20119 27285 20131 27319
rect 20073 27279 20131 27285
rect 20806 27276 20812 27328
rect 20864 27316 20870 27328
rect 22547 27316 22575 27344
rect 22922 27316 22928 27328
rect 20864 27288 22928 27316
rect 20864 27276 20870 27288
rect 22922 27276 22928 27288
rect 22980 27316 22986 27328
rect 23609 27316 23637 27347
rect 23750 27344 23756 27356
rect 23808 27344 23814 27396
rect 24596 27384 24624 27415
rect 24670 27412 24676 27464
rect 24728 27452 24734 27464
rect 24949 27455 25007 27461
rect 24949 27452 24961 27455
rect 24728 27424 24961 27452
rect 24728 27412 24734 27424
rect 24949 27421 24961 27424
rect 24995 27421 25007 27455
rect 25409 27455 25467 27461
rect 25409 27452 25421 27455
rect 24949 27415 25007 27421
rect 25332 27424 25421 27452
rect 25332 27384 25360 27424
rect 25409 27421 25421 27424
rect 25455 27421 25467 27455
rect 25409 27415 25467 27421
rect 25498 27412 25504 27464
rect 25556 27452 25562 27464
rect 25774 27452 25780 27464
rect 25556 27424 25780 27452
rect 25556 27412 25562 27424
rect 25774 27412 25780 27424
rect 25832 27412 25838 27464
rect 25958 27412 25964 27464
rect 26016 27412 26022 27464
rect 26068 27461 26096 27492
rect 26326 27480 26332 27532
rect 26384 27480 26390 27532
rect 26528 27461 26556 27560
rect 26620 27492 27108 27520
rect 26053 27455 26111 27461
rect 26053 27421 26065 27455
rect 26099 27421 26111 27455
rect 26053 27415 26111 27421
rect 26513 27455 26571 27461
rect 26513 27421 26525 27455
rect 26559 27421 26571 27455
rect 26513 27415 26571 27421
rect 25976 27384 26004 27412
rect 24596 27356 25360 27384
rect 22980 27288 23637 27316
rect 25332 27316 25360 27356
rect 25792 27356 26004 27384
rect 25792 27328 25820 27356
rect 26234 27344 26240 27396
rect 26292 27384 26298 27396
rect 26620 27384 26648 27492
rect 26786 27412 26792 27464
rect 26844 27412 26850 27464
rect 27080 27461 27108 27492
rect 26973 27455 27031 27461
rect 26973 27421 26985 27455
rect 27019 27421 27031 27455
rect 26973 27415 27031 27421
rect 27065 27455 27123 27461
rect 27065 27421 27077 27455
rect 27111 27421 27123 27455
rect 27065 27415 27123 27421
rect 27249 27455 27307 27461
rect 27249 27421 27261 27455
rect 27295 27421 27307 27455
rect 27249 27415 27307 27421
rect 26988 27384 27016 27415
rect 27264 27384 27292 27415
rect 26292 27356 26648 27384
rect 26712 27356 27292 27384
rect 26292 27344 26298 27356
rect 25774 27316 25780 27328
rect 25332 27288 25780 27316
rect 22980 27276 22986 27288
rect 25774 27276 25780 27288
rect 25832 27276 25838 27328
rect 25958 27276 25964 27328
rect 26016 27276 26022 27328
rect 26712 27325 26740 27356
rect 26697 27319 26755 27325
rect 26697 27285 26709 27319
rect 26743 27285 26755 27319
rect 26697 27279 26755 27285
rect 1104 27226 28152 27248
rect 1104 27174 4874 27226
rect 4926 27174 4938 27226
rect 4990 27174 5002 27226
rect 5054 27174 5066 27226
rect 5118 27174 5130 27226
rect 5182 27174 28152 27226
rect 1104 27152 28152 27174
rect 5077 27115 5135 27121
rect 5077 27081 5089 27115
rect 5123 27112 5135 27115
rect 5258 27112 5264 27124
rect 5123 27084 5264 27112
rect 5123 27081 5135 27084
rect 5077 27075 5135 27081
rect 5258 27072 5264 27084
rect 5316 27112 5322 27124
rect 5971 27115 6029 27121
rect 5971 27112 5983 27115
rect 5316 27084 5983 27112
rect 5316 27072 5322 27084
rect 5971 27081 5983 27084
rect 6017 27081 6029 27115
rect 11054 27112 11060 27124
rect 5971 27075 6029 27081
rect 10888 27084 11060 27112
rect 2774 27004 2780 27056
rect 2832 27004 2838 27056
rect 2977 27047 3035 27053
rect 2977 27044 2989 27047
rect 2884 27016 2989 27044
rect 2038 26936 2044 26988
rect 2096 26976 2102 26988
rect 2225 26979 2283 26985
rect 2225 26976 2237 26979
rect 2096 26948 2237 26976
rect 2096 26936 2102 26948
rect 2225 26945 2237 26948
rect 2271 26945 2283 26979
rect 2884 26976 2912 27016
rect 2977 27013 2989 27016
rect 3023 27013 3035 27047
rect 5442 27044 5448 27056
rect 2977 27007 3035 27013
rect 3988 27016 5448 27044
rect 2225 26939 2283 26945
rect 2608 26948 2912 26976
rect 2608 26920 2636 26948
rect 3510 26936 3516 26988
rect 3568 26936 3574 26988
rect 3988 26985 4016 27016
rect 5442 27004 5448 27016
rect 5500 27004 5506 27056
rect 6181 27047 6239 27053
rect 6181 27013 6193 27047
rect 6227 27044 6239 27047
rect 6638 27044 6644 27056
rect 6227 27016 6644 27044
rect 6227 27013 6239 27016
rect 6181 27007 6239 27013
rect 6638 27004 6644 27016
rect 6696 27004 6702 27056
rect 7650 27044 7656 27056
rect 6748 27016 7656 27044
rect 3697 26979 3755 26985
rect 3697 26945 3709 26979
rect 3743 26976 3755 26979
rect 3973 26979 4031 26985
rect 3973 26976 3985 26979
rect 3743 26948 3985 26976
rect 3743 26945 3755 26948
rect 3697 26939 3755 26945
rect 3973 26945 3985 26948
rect 4019 26945 4031 26979
rect 3973 26939 4031 26945
rect 4709 26979 4767 26985
rect 4709 26945 4721 26979
rect 4755 26976 4767 26979
rect 5353 26979 5411 26985
rect 5353 26976 5365 26979
rect 4755 26948 5365 26976
rect 4755 26945 4767 26948
rect 4709 26939 4767 26945
rect 5353 26945 5365 26948
rect 5399 26945 5411 26979
rect 5353 26939 5411 26945
rect 2130 26868 2136 26920
rect 2188 26868 2194 26920
rect 2590 26868 2596 26920
rect 2648 26868 2654 26920
rect 3237 26911 3295 26917
rect 3237 26908 3249 26911
rect 3160 26880 3249 26908
rect 2148 26840 2176 26868
rect 3050 26840 3056 26852
rect 2148 26812 3056 26840
rect 3050 26800 3056 26812
rect 3108 26800 3114 26852
rect 2498 26732 2504 26784
rect 2556 26772 2562 26784
rect 3160 26781 3188 26880
rect 3237 26877 3249 26880
rect 3283 26908 3295 26911
rect 3786 26908 3792 26920
rect 3283 26880 3792 26908
rect 3283 26877 3295 26880
rect 3237 26871 3295 26877
rect 3786 26868 3792 26880
rect 3844 26868 3850 26920
rect 3878 26868 3884 26920
rect 3936 26868 3942 26920
rect 3513 26843 3571 26849
rect 3513 26809 3525 26843
rect 3559 26840 3571 26843
rect 4724 26840 4752 26939
rect 5534 26936 5540 26988
rect 5592 26936 5598 26988
rect 6546 26936 6552 26988
rect 6604 26976 6610 26988
rect 6748 26976 6776 27016
rect 6604 26948 6776 26976
rect 6604 26936 6610 26948
rect 6914 26936 6920 26988
rect 6972 26976 6978 26988
rect 7392 26985 7420 27016
rect 7650 27004 7656 27016
rect 7708 27044 7714 27056
rect 10888 27044 10916 27084
rect 11054 27072 11060 27084
rect 11112 27072 11118 27124
rect 11241 27115 11299 27121
rect 11241 27081 11253 27115
rect 11287 27112 11299 27115
rect 11287 27084 12204 27112
rect 11287 27081 11299 27084
rect 11241 27075 11299 27081
rect 11900 27053 11928 27084
rect 11669 27047 11727 27053
rect 11669 27044 11681 27047
rect 7708 27016 10916 27044
rect 10980 27016 11681 27044
rect 7708 27004 7714 27016
rect 10980 26988 11008 27016
rect 11669 27013 11681 27016
rect 11715 27013 11727 27047
rect 11669 27007 11727 27013
rect 11885 27047 11943 27053
rect 11885 27013 11897 27047
rect 11931 27013 11943 27047
rect 11885 27007 11943 27013
rect 11974 27004 11980 27056
rect 12032 27004 12038 27056
rect 12176 27053 12204 27084
rect 12342 27072 12348 27124
rect 12400 27112 12406 27124
rect 12529 27115 12587 27121
rect 12529 27112 12541 27115
rect 12400 27084 12541 27112
rect 12400 27072 12406 27084
rect 12529 27081 12541 27084
rect 12575 27081 12587 27115
rect 12529 27075 12587 27081
rect 17402 27072 17408 27124
rect 17460 27072 17466 27124
rect 18046 27072 18052 27124
rect 18104 27072 18110 27124
rect 18138 27072 18144 27124
rect 18196 27072 18202 27124
rect 18693 27115 18751 27121
rect 18432 27084 18644 27112
rect 12161 27047 12219 27053
rect 12161 27013 12173 27047
rect 12207 27013 12219 27047
rect 12986 27044 12992 27056
rect 12161 27007 12219 27013
rect 12268 27016 12992 27044
rect 7009 26979 7067 26985
rect 7009 26976 7021 26979
rect 6972 26948 7021 26976
rect 6972 26936 6978 26948
rect 7009 26945 7021 26948
rect 7055 26976 7067 26979
rect 7101 26979 7159 26985
rect 7101 26976 7113 26979
rect 7055 26948 7113 26976
rect 7055 26945 7067 26948
rect 7009 26939 7067 26945
rect 7101 26945 7113 26948
rect 7147 26945 7159 26979
rect 7101 26939 7159 26945
rect 7377 26979 7435 26985
rect 7377 26945 7389 26979
rect 7423 26945 7435 26979
rect 7377 26939 7435 26945
rect 9122 26936 9128 26988
rect 9180 26936 9186 26988
rect 10594 26936 10600 26988
rect 10652 26976 10658 26988
rect 10689 26979 10747 26985
rect 10689 26976 10701 26979
rect 10652 26948 10701 26976
rect 10652 26936 10658 26948
rect 10689 26945 10701 26948
rect 10735 26945 10747 26979
rect 10689 26939 10747 26945
rect 10778 26936 10784 26988
rect 10836 26936 10842 26988
rect 10962 26936 10968 26988
rect 11020 26936 11026 26988
rect 11054 26936 11060 26988
rect 11112 26976 11118 26988
rect 11149 26979 11207 26985
rect 11149 26976 11161 26979
rect 11112 26948 11161 26976
rect 11112 26936 11118 26948
rect 11149 26945 11161 26948
rect 11195 26976 11207 26979
rect 12268 26976 12296 27016
rect 12986 27004 12992 27016
rect 13044 27004 13050 27056
rect 16942 27004 16948 27056
rect 17000 27044 17006 27056
rect 18064 27044 18092 27072
rect 18293 27047 18351 27053
rect 18293 27044 18305 27047
rect 17000 27016 17908 27044
rect 18064 27016 18305 27044
rect 17000 27004 17006 27016
rect 11195 26948 12296 26976
rect 12345 26979 12403 26985
rect 11195 26945 11207 26948
rect 11149 26939 11207 26945
rect 12345 26945 12357 26979
rect 12391 26976 12403 26979
rect 12437 26979 12495 26985
rect 12437 26976 12449 26979
rect 12391 26948 12449 26976
rect 12391 26945 12403 26948
rect 12345 26939 12403 26945
rect 12437 26945 12449 26948
rect 12483 26945 12495 26979
rect 12437 26939 12495 26945
rect 12710 26936 12716 26988
rect 12768 26936 12774 26988
rect 17328 26985 17356 27016
rect 17880 26985 17908 27016
rect 18293 27013 18305 27016
rect 18339 27013 18351 27047
rect 18293 27007 18351 27013
rect 17313 26979 17371 26985
rect 17313 26945 17325 26979
rect 17359 26945 17371 26979
rect 17313 26939 17371 26945
rect 17497 26979 17555 26985
rect 17497 26945 17509 26979
rect 17543 26945 17555 26979
rect 17497 26939 17555 26945
rect 17865 26979 17923 26985
rect 17865 26945 17877 26979
rect 17911 26976 17923 26979
rect 17954 26976 17960 26988
rect 17911 26948 17960 26976
rect 17911 26945 17923 26948
rect 17865 26939 17923 26945
rect 4798 26868 4804 26920
rect 4856 26868 4862 26920
rect 5261 26911 5319 26917
rect 5261 26877 5273 26911
rect 5307 26877 5319 26911
rect 5261 26871 5319 26877
rect 3559 26812 4752 26840
rect 5276 26840 5304 26871
rect 5442 26868 5448 26920
rect 5500 26868 5506 26920
rect 5718 26868 5724 26920
rect 5776 26868 5782 26920
rect 6822 26868 6828 26920
rect 6880 26908 6886 26920
rect 7193 26911 7251 26917
rect 7193 26908 7205 26911
rect 6880 26880 7205 26908
rect 6880 26868 6886 26880
rect 7193 26877 7205 26880
rect 7239 26877 7251 26911
rect 7193 26871 7251 26877
rect 9217 26911 9275 26917
rect 9217 26877 9229 26911
rect 9263 26908 9275 26911
rect 9769 26911 9827 26917
rect 9769 26908 9781 26911
rect 9263 26880 9781 26908
rect 9263 26877 9275 26880
rect 9217 26871 9275 26877
rect 9769 26877 9781 26880
rect 9815 26877 9827 26911
rect 9769 26871 9827 26877
rect 5810 26840 5816 26852
rect 5276 26812 5816 26840
rect 3559 26809 3571 26812
rect 3513 26803 3571 26809
rect 5810 26800 5816 26812
rect 5868 26800 5874 26852
rect 5902 26800 5908 26852
rect 5960 26840 5966 26852
rect 6687 26843 6745 26849
rect 6687 26840 6699 26843
rect 5960 26812 6699 26840
rect 5960 26800 5966 26812
rect 6687 26809 6699 26812
rect 6733 26840 6745 26843
rect 7006 26840 7012 26852
rect 6733 26812 7012 26840
rect 6733 26809 6745 26812
rect 6687 26803 6745 26809
rect 7006 26800 7012 26812
rect 7064 26840 7070 26852
rect 9784 26840 9812 26871
rect 9858 26868 9864 26920
rect 9916 26868 9922 26920
rect 10229 26911 10287 26917
rect 10229 26877 10241 26911
rect 10275 26877 10287 26911
rect 10229 26871 10287 26877
rect 10873 26911 10931 26917
rect 10873 26877 10885 26911
rect 10919 26877 10931 26911
rect 17512 26908 17540 26939
rect 17954 26936 17960 26948
rect 18012 26936 18018 26988
rect 18049 26979 18107 26985
rect 18049 26945 18061 26979
rect 18095 26976 18107 26979
rect 18432 26976 18460 27084
rect 18506 27004 18512 27056
rect 18564 27004 18570 27056
rect 18616 27044 18644 27084
rect 18693 27081 18705 27115
rect 18739 27112 18751 27115
rect 19426 27112 19432 27124
rect 18739 27084 19432 27112
rect 18739 27081 18751 27084
rect 18693 27075 18751 27081
rect 19426 27072 19432 27084
rect 19484 27072 19490 27124
rect 19613 27115 19671 27121
rect 19613 27081 19625 27115
rect 19659 27112 19671 27115
rect 20346 27112 20352 27124
rect 19659 27084 20352 27112
rect 19659 27081 19671 27084
rect 19613 27075 19671 27081
rect 19628 27044 19656 27075
rect 20346 27072 20352 27084
rect 20404 27072 20410 27124
rect 20990 27072 20996 27124
rect 21048 27072 21054 27124
rect 21542 27072 21548 27124
rect 21600 27112 21606 27124
rect 22189 27115 22247 27121
rect 22189 27112 22201 27115
rect 21600 27084 22201 27112
rect 21600 27072 21606 27084
rect 22189 27081 22201 27084
rect 22235 27081 22247 27115
rect 22189 27075 22247 27081
rect 22373 27115 22431 27121
rect 22373 27081 22385 27115
rect 22419 27112 22431 27115
rect 22646 27112 22652 27124
rect 22419 27084 22652 27112
rect 22419 27081 22431 27084
rect 22373 27075 22431 27081
rect 22646 27072 22652 27084
rect 22704 27072 22710 27124
rect 23201 27115 23259 27121
rect 23201 27081 23213 27115
rect 23247 27112 23259 27115
rect 23290 27112 23296 27124
rect 23247 27084 23296 27112
rect 23247 27081 23259 27084
rect 23201 27075 23259 27081
rect 23290 27072 23296 27084
rect 23348 27072 23354 27124
rect 24210 27072 24216 27124
rect 24268 27112 24274 27124
rect 24762 27112 24768 27124
rect 24268 27084 24768 27112
rect 24268 27072 24274 27084
rect 24762 27072 24768 27084
rect 24820 27072 24826 27124
rect 24949 27115 25007 27121
rect 24949 27081 24961 27115
rect 24995 27112 25007 27115
rect 25866 27112 25872 27124
rect 24995 27084 25872 27112
rect 24995 27081 25007 27084
rect 24949 27075 25007 27081
rect 25866 27072 25872 27084
rect 25924 27072 25930 27124
rect 25961 27115 26019 27121
rect 25961 27081 25973 27115
rect 26007 27112 26019 27115
rect 26050 27112 26056 27124
rect 26007 27084 26056 27112
rect 26007 27081 26019 27084
rect 25961 27075 26019 27081
rect 26050 27072 26056 27084
rect 26108 27072 26114 27124
rect 19978 27044 19984 27056
rect 18616 27016 19656 27044
rect 19720 27016 19984 27044
rect 18095 26948 18460 26976
rect 18601 26979 18659 26985
rect 18095 26945 18107 26948
rect 18049 26939 18107 26945
rect 18601 26945 18613 26979
rect 18647 26945 18659 26979
rect 18601 26939 18659 26945
rect 18616 26908 18644 26939
rect 18690 26936 18696 26988
rect 18748 26976 18754 26988
rect 18785 26979 18843 26985
rect 18785 26976 18797 26979
rect 18748 26948 18797 26976
rect 18748 26936 18754 26948
rect 18785 26945 18797 26948
rect 18831 26945 18843 26979
rect 18785 26939 18843 26945
rect 19061 26979 19119 26985
rect 19061 26945 19073 26979
rect 19107 26976 19119 26979
rect 19107 26948 19334 26976
rect 19107 26945 19119 26948
rect 19061 26939 19119 26945
rect 19153 26911 19211 26917
rect 17512 26880 18920 26908
rect 10873 26871 10931 26877
rect 9950 26840 9956 26852
rect 7064 26812 7144 26840
rect 9784 26812 9956 26840
rect 7064 26800 7070 26812
rect 2961 26775 3019 26781
rect 2961 26772 2973 26775
rect 2556 26744 2973 26772
rect 2556 26732 2562 26744
rect 2961 26741 2973 26744
rect 3007 26741 3019 26775
rect 2961 26735 3019 26741
rect 3145 26775 3203 26781
rect 3145 26741 3157 26775
rect 3191 26741 3203 26775
rect 3145 26735 3203 26741
rect 4249 26775 4307 26781
rect 4249 26741 4261 26775
rect 4295 26772 4307 26775
rect 4706 26772 4712 26784
rect 4295 26744 4712 26772
rect 4295 26741 4307 26744
rect 4249 26735 4307 26741
rect 4706 26732 4712 26744
rect 4764 26732 4770 26784
rect 4982 26732 4988 26784
rect 5040 26772 5046 26784
rect 5626 26772 5632 26784
rect 5040 26744 5632 26772
rect 5040 26732 5046 26744
rect 5626 26732 5632 26744
rect 5684 26772 5690 26784
rect 5997 26775 6055 26781
rect 5997 26772 6009 26775
rect 5684 26744 6009 26772
rect 5684 26732 5690 26744
rect 5997 26741 6009 26744
rect 6043 26741 6055 26775
rect 5997 26735 6055 26741
rect 6178 26732 6184 26784
rect 6236 26772 6242 26784
rect 6822 26772 6828 26784
rect 6236 26744 6828 26772
rect 6236 26732 6242 26744
rect 6822 26732 6828 26744
rect 6880 26732 6886 26784
rect 6914 26732 6920 26784
rect 6972 26732 6978 26784
rect 7116 26781 7144 26812
rect 9950 26800 9956 26812
rect 10008 26800 10014 26852
rect 10244 26840 10272 26871
rect 10410 26840 10416 26852
rect 10244 26812 10416 26840
rect 10410 26800 10416 26812
rect 10468 26840 10474 26852
rect 10468 26812 10640 26840
rect 10468 26800 10474 26812
rect 10612 26784 10640 26812
rect 7101 26775 7159 26781
rect 7101 26741 7113 26775
rect 7147 26741 7159 26775
rect 7101 26735 7159 26741
rect 7561 26775 7619 26781
rect 7561 26741 7573 26775
rect 7607 26772 7619 26775
rect 7650 26772 7656 26784
rect 7607 26744 7656 26772
rect 7607 26741 7619 26744
rect 7561 26735 7619 26741
rect 7650 26732 7656 26744
rect 7708 26732 7714 26784
rect 8754 26732 8760 26784
rect 8812 26772 8818 26784
rect 8849 26775 8907 26781
rect 8849 26772 8861 26775
rect 8812 26744 8861 26772
rect 8812 26732 8818 26744
rect 8849 26741 8861 26744
rect 8895 26741 8907 26775
rect 8849 26735 8907 26741
rect 9585 26775 9643 26781
rect 9585 26741 9597 26775
rect 9631 26772 9643 26775
rect 9766 26772 9772 26784
rect 9631 26744 9772 26772
rect 9631 26741 9643 26744
rect 9585 26735 9643 26741
rect 9766 26732 9772 26744
rect 9824 26732 9830 26784
rect 10226 26732 10232 26784
rect 10284 26772 10290 26784
rect 10505 26775 10563 26781
rect 10505 26772 10517 26775
rect 10284 26744 10517 26772
rect 10284 26732 10290 26744
rect 10505 26741 10517 26744
rect 10551 26741 10563 26775
rect 10505 26735 10563 26741
rect 10594 26732 10600 26784
rect 10652 26732 10658 26784
rect 10888 26772 10916 26871
rect 17862 26800 17868 26852
rect 17920 26800 17926 26852
rect 17954 26800 17960 26852
rect 18012 26840 18018 26852
rect 18782 26840 18788 26852
rect 18012 26812 18788 26840
rect 18012 26800 18018 26812
rect 18782 26800 18788 26812
rect 18840 26800 18846 26852
rect 18892 26849 18920 26880
rect 19153 26877 19165 26911
rect 19199 26877 19211 26911
rect 19306 26908 19334 26948
rect 19518 26936 19524 26988
rect 19576 26976 19582 26988
rect 19720 26976 19748 27016
rect 19978 27004 19984 27016
rect 20036 27004 20042 27056
rect 20898 27044 20904 27056
rect 20364 27016 20904 27044
rect 19576 26948 19748 26976
rect 19576 26936 19582 26948
rect 19794 26936 19800 26988
rect 19852 26976 19858 26988
rect 19852 26948 20208 26976
rect 19852 26936 19858 26948
rect 19812 26908 19840 26936
rect 19306 26880 19840 26908
rect 19153 26871 19211 26877
rect 18877 26843 18935 26849
rect 18877 26809 18889 26843
rect 18923 26809 18935 26843
rect 18877 26803 18935 26809
rect 11238 26772 11244 26784
rect 10888 26744 11244 26772
rect 11238 26732 11244 26744
rect 11296 26732 11302 26784
rect 11514 26732 11520 26784
rect 11572 26732 11578 26784
rect 11698 26732 11704 26784
rect 11756 26732 11762 26784
rect 12526 26732 12532 26784
rect 12584 26772 12590 26784
rect 12713 26775 12771 26781
rect 12713 26772 12725 26775
rect 12584 26744 12725 26772
rect 12584 26732 12590 26744
rect 12713 26741 12725 26744
rect 12759 26741 12771 26775
rect 12713 26735 12771 26741
rect 18322 26732 18328 26784
rect 18380 26732 18386 26784
rect 18506 26732 18512 26784
rect 18564 26772 18570 26784
rect 19061 26775 19119 26781
rect 19061 26772 19073 26775
rect 18564 26744 19073 26772
rect 18564 26732 18570 26744
rect 19061 26741 19073 26744
rect 19107 26741 19119 26775
rect 19168 26772 19196 26871
rect 19978 26868 19984 26920
rect 20036 26868 20042 26920
rect 20180 26908 20208 26948
rect 20254 26936 20260 26988
rect 20312 26936 20318 26988
rect 20364 26985 20392 27016
rect 20898 27004 20904 27016
rect 20956 27044 20962 27056
rect 21085 27047 21143 27053
rect 21085 27044 21097 27047
rect 20956 27016 21097 27044
rect 20956 27004 20962 27016
rect 21085 27013 21097 27016
rect 21131 27013 21143 27047
rect 21910 27044 21916 27056
rect 21085 27007 21143 27013
rect 21314 27016 21916 27044
rect 20349 26979 20407 26985
rect 20349 26945 20361 26979
rect 20395 26945 20407 26979
rect 20349 26939 20407 26945
rect 20533 26979 20591 26985
rect 20533 26945 20545 26979
rect 20579 26945 20591 26979
rect 20533 26939 20591 26945
rect 20438 26908 20444 26920
rect 20180 26880 20444 26908
rect 20438 26868 20444 26880
rect 20496 26868 20502 26920
rect 19242 26800 19248 26852
rect 19300 26840 19306 26852
rect 20548 26840 20576 26939
rect 20622 26936 20628 26988
rect 20680 26976 20686 26988
rect 20809 26979 20867 26985
rect 20809 26976 20821 26979
rect 20680 26948 20821 26976
rect 20680 26936 20686 26948
rect 20809 26945 20821 26948
rect 20855 26976 20867 26979
rect 20990 26976 20996 26988
rect 20855 26948 20996 26976
rect 20855 26945 20867 26948
rect 20809 26939 20867 26945
rect 20990 26936 20996 26948
rect 21048 26976 21054 26988
rect 21314 26985 21342 27016
rect 21910 27004 21916 27016
rect 21968 27004 21974 27056
rect 22005 27047 22063 27053
rect 22005 27013 22017 27047
rect 22051 27044 22063 27047
rect 22278 27044 22284 27056
rect 22051 27016 22284 27044
rect 22051 27013 22063 27016
rect 22005 27007 22063 27013
rect 22278 27004 22284 27016
rect 22336 27004 22342 27056
rect 22462 27004 22468 27056
rect 22520 27044 22526 27056
rect 23106 27044 23112 27056
rect 22520 27016 23112 27044
rect 22520 27004 22526 27016
rect 23106 27004 23112 27016
rect 23164 27004 23170 27056
rect 25406 27004 25412 27056
rect 25464 27004 25470 27056
rect 26786 27044 26792 27056
rect 25884 27016 26792 27044
rect 25884 26988 25912 27016
rect 26786 27004 26792 27016
rect 26844 27004 26850 27056
rect 21299 26979 21357 26985
rect 21299 26976 21311 26979
rect 21048 26948 21311 26976
rect 21048 26936 21054 26948
rect 21299 26945 21311 26948
rect 21345 26945 21357 26979
rect 21299 26939 21357 26945
rect 21450 26936 21456 26988
rect 21508 26936 21514 26988
rect 22097 26979 22155 26985
rect 22097 26945 22109 26979
rect 22143 26945 22155 26979
rect 22097 26939 22155 26945
rect 20717 26911 20775 26917
rect 20717 26877 20729 26911
rect 20763 26908 20775 26911
rect 22112 26908 22140 26939
rect 22646 26936 22652 26988
rect 22704 26936 22710 26988
rect 22922 26936 22928 26988
rect 22980 26936 22986 26988
rect 23014 26936 23020 26988
rect 23072 26976 23078 26988
rect 23072 26948 23244 26976
rect 23072 26936 23078 26948
rect 22557 26911 22615 26917
rect 22557 26908 22569 26911
rect 20763 26880 22569 26908
rect 20763 26877 20775 26880
rect 20717 26871 20775 26877
rect 22557 26877 22569 26880
rect 22603 26877 22615 26911
rect 22557 26871 22615 26877
rect 19300 26812 20576 26840
rect 19300 26800 19306 26812
rect 20622 26800 20628 26852
rect 20680 26800 20686 26852
rect 21818 26840 21824 26852
rect 20732 26812 21824 26840
rect 20162 26772 20168 26784
rect 19168 26744 20168 26772
rect 19061 26735 19119 26741
rect 20162 26732 20168 26744
rect 20220 26732 20226 26784
rect 20438 26732 20444 26784
rect 20496 26772 20502 26784
rect 20732 26772 20760 26812
rect 21818 26800 21824 26812
rect 21876 26800 21882 26852
rect 22278 26800 22284 26852
rect 22336 26840 22342 26852
rect 23216 26840 23244 26948
rect 23658 26936 23664 26988
rect 23716 26976 23722 26988
rect 24121 26979 24179 26985
rect 24121 26976 24133 26979
rect 23716 26948 24133 26976
rect 23716 26936 23722 26948
rect 24121 26945 24133 26948
rect 24167 26976 24179 26979
rect 24394 26976 24400 26988
rect 24167 26948 24400 26976
rect 24167 26945 24179 26948
rect 24121 26939 24179 26945
rect 24394 26936 24400 26948
rect 24452 26936 24458 26988
rect 24581 26979 24639 26985
rect 24581 26945 24593 26979
rect 24627 26976 24639 26979
rect 24670 26976 24676 26988
rect 24627 26948 24676 26976
rect 24627 26945 24639 26948
rect 24581 26939 24639 26945
rect 24670 26936 24676 26948
rect 24728 26936 24734 26988
rect 24762 26936 24768 26988
rect 24820 26976 24826 26988
rect 24857 26979 24915 26985
rect 24857 26976 24869 26979
rect 24820 26948 24869 26976
rect 24820 26936 24826 26948
rect 24857 26945 24869 26948
rect 24903 26945 24915 26979
rect 24857 26939 24915 26945
rect 24946 26936 24952 26988
rect 25004 26976 25010 26988
rect 25041 26979 25099 26985
rect 25041 26976 25053 26979
rect 25004 26948 25053 26976
rect 25004 26936 25010 26948
rect 25041 26945 25053 26948
rect 25087 26945 25099 26979
rect 25041 26939 25099 26945
rect 25130 26936 25136 26988
rect 25188 26976 25194 26988
rect 25317 26979 25375 26985
rect 25317 26976 25329 26979
rect 25188 26948 25329 26976
rect 25188 26936 25194 26948
rect 25317 26945 25329 26948
rect 25363 26945 25375 26979
rect 25317 26939 25375 26945
rect 25501 26979 25559 26985
rect 25501 26945 25513 26979
rect 25547 26976 25559 26979
rect 25547 26948 25636 26976
rect 25547 26945 25559 26948
rect 25501 26939 25559 26945
rect 24486 26868 24492 26920
rect 24544 26908 24550 26920
rect 25222 26908 25228 26920
rect 24544 26880 25228 26908
rect 24544 26868 24550 26880
rect 25222 26868 25228 26880
rect 25280 26868 25286 26920
rect 25608 26908 25636 26948
rect 25866 26936 25872 26988
rect 25924 26936 25930 26988
rect 25958 26936 25964 26988
rect 26016 26976 26022 26988
rect 26053 26979 26111 26985
rect 26053 26976 26065 26979
rect 26016 26948 26065 26976
rect 26016 26936 26022 26948
rect 26053 26945 26065 26948
rect 26099 26976 26111 26979
rect 26145 26979 26203 26985
rect 26145 26976 26157 26979
rect 26099 26948 26157 26976
rect 26099 26945 26111 26948
rect 26053 26939 26111 26945
rect 26145 26945 26157 26948
rect 26191 26945 26203 26979
rect 26145 26939 26203 26945
rect 26234 26936 26240 26988
rect 26292 26976 26298 26988
rect 26329 26979 26387 26985
rect 26329 26976 26341 26979
rect 26292 26948 26341 26976
rect 26292 26936 26298 26948
rect 26329 26945 26341 26948
rect 26375 26945 26387 26979
rect 26329 26939 26387 26945
rect 26252 26908 26280 26936
rect 25608 26880 26280 26908
rect 25590 26840 25596 26852
rect 22336 26812 25596 26840
rect 22336 26800 22342 26812
rect 25590 26800 25596 26812
rect 25648 26800 25654 26852
rect 26142 26800 26148 26852
rect 26200 26800 26206 26852
rect 20496 26744 20760 26772
rect 20496 26732 20502 26744
rect 24210 26732 24216 26784
rect 24268 26732 24274 26784
rect 1104 26682 28152 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 28152 26682
rect 1104 26608 28152 26630
rect 3050 26528 3056 26580
rect 3108 26568 3114 26580
rect 3108 26540 3648 26568
rect 3108 26528 3114 26540
rect 2130 26500 2136 26512
rect 1780 26472 2136 26500
rect 1780 26373 1808 26472
rect 2130 26460 2136 26472
rect 2188 26460 2194 26512
rect 2590 26460 2596 26512
rect 2648 26500 2654 26512
rect 3145 26503 3203 26509
rect 2648 26472 3096 26500
rect 2648 26460 2654 26472
rect 3068 26432 3096 26472
rect 3145 26469 3157 26503
rect 3191 26500 3203 26503
rect 3510 26500 3516 26512
rect 3191 26472 3516 26500
rect 3191 26469 3203 26472
rect 3145 26463 3203 26469
rect 3510 26460 3516 26472
rect 3568 26460 3574 26512
rect 1964 26404 3020 26432
rect 3068 26404 3188 26432
rect 1765 26367 1823 26373
rect 1765 26333 1777 26367
rect 1811 26333 1823 26367
rect 1964 26366 1992 26404
rect 1765 26327 1823 26333
rect 1872 26338 1992 26366
rect 2869 26367 2927 26373
rect 2869 26364 2881 26367
rect 1872 26296 1900 26338
rect 2746 26336 2881 26364
rect 1780 26268 1900 26296
rect 1780 26240 1808 26268
rect 2498 26256 2504 26308
rect 2556 26296 2562 26308
rect 2746 26296 2774 26336
rect 2869 26333 2881 26336
rect 2915 26333 2927 26367
rect 2869 26327 2927 26333
rect 2556 26268 2774 26296
rect 2992 26296 3020 26404
rect 3160 26373 3188 26404
rect 3145 26367 3203 26373
rect 3145 26333 3157 26367
rect 3191 26333 3203 26367
rect 3528 26364 3556 26460
rect 3620 26432 3648 26540
rect 3878 26528 3884 26580
rect 3936 26568 3942 26580
rect 3973 26571 4031 26577
rect 3973 26568 3985 26571
rect 3936 26540 3985 26568
rect 3936 26528 3942 26540
rect 3973 26537 3985 26540
rect 4019 26537 4031 26571
rect 3973 26531 4031 26537
rect 4798 26528 4804 26580
rect 4856 26568 4862 26580
rect 5445 26571 5503 26577
rect 5445 26568 5457 26571
rect 4856 26540 5457 26568
rect 4856 26528 4862 26540
rect 5445 26537 5457 26540
rect 5491 26537 5503 26571
rect 5445 26531 5503 26537
rect 7006 26528 7012 26580
rect 7064 26528 7070 26580
rect 9858 26568 9864 26580
rect 7576 26540 9864 26568
rect 4062 26460 4068 26512
rect 4120 26500 4126 26512
rect 6546 26500 6552 26512
rect 4120 26472 6552 26500
rect 4120 26460 4126 26472
rect 4614 26432 4620 26444
rect 3620 26404 4620 26432
rect 4614 26392 4620 26404
rect 4672 26432 4678 26444
rect 4672 26404 5120 26432
rect 4672 26392 4678 26404
rect 3789 26367 3847 26373
rect 3789 26364 3801 26367
rect 3528 26336 3801 26364
rect 3145 26327 3203 26333
rect 3789 26333 3801 26336
rect 3835 26333 3847 26367
rect 3789 26327 3847 26333
rect 3878 26324 3884 26376
rect 3936 26364 3942 26376
rect 3973 26367 4031 26373
rect 3973 26364 3985 26367
rect 3936 26336 3985 26364
rect 3936 26324 3942 26336
rect 3973 26333 3985 26336
rect 4019 26333 4031 26367
rect 3973 26327 4031 26333
rect 4982 26324 4988 26376
rect 5040 26324 5046 26376
rect 4798 26296 4804 26308
rect 2992 26268 4804 26296
rect 2556 26256 2562 26268
rect 4798 26256 4804 26268
rect 4856 26296 4862 26308
rect 5000 26296 5028 26324
rect 5092 26305 5120 26404
rect 5166 26392 5172 26444
rect 5224 26432 5230 26444
rect 5224 26404 5672 26432
rect 5224 26392 5230 26404
rect 5258 26324 5264 26376
rect 5316 26324 5322 26376
rect 5350 26324 5356 26376
rect 5408 26324 5414 26376
rect 5534 26324 5540 26376
rect 5592 26324 5598 26376
rect 5644 26373 5672 26404
rect 5629 26367 5687 26373
rect 5629 26333 5641 26367
rect 5675 26333 5687 26367
rect 5629 26327 5687 26333
rect 5810 26324 5816 26376
rect 5868 26324 5874 26376
rect 6104 26364 6132 26472
rect 6546 26460 6552 26472
rect 6604 26460 6610 26512
rect 6638 26460 6644 26512
rect 6696 26500 6702 26512
rect 6696 26472 6868 26500
rect 6696 26460 6702 26472
rect 6273 26435 6331 26441
rect 6273 26401 6285 26435
rect 6319 26432 6331 26435
rect 6733 26435 6791 26441
rect 6733 26432 6745 26435
rect 6319 26404 6745 26432
rect 6319 26401 6331 26404
rect 6273 26395 6331 26401
rect 6733 26401 6745 26404
rect 6779 26401 6791 26435
rect 6733 26395 6791 26401
rect 6181 26367 6239 26373
rect 6181 26364 6193 26367
rect 6104 26336 6193 26364
rect 6181 26333 6193 26336
rect 6227 26333 6239 26367
rect 6181 26327 6239 26333
rect 6638 26324 6644 26376
rect 6696 26324 6702 26376
rect 6840 26373 6868 26472
rect 6914 26392 6920 26444
rect 6972 26432 6978 26444
rect 6972 26404 7512 26432
rect 6972 26392 6978 26404
rect 7484 26373 7512 26404
rect 6825 26367 6883 26373
rect 6825 26333 6837 26367
rect 6871 26364 6883 26367
rect 7101 26367 7159 26373
rect 7101 26364 7113 26367
rect 6871 26336 7113 26364
rect 6871 26333 6883 26336
rect 6825 26327 6883 26333
rect 7101 26333 7113 26336
rect 7147 26333 7159 26367
rect 7101 26327 7159 26333
rect 7469 26367 7527 26373
rect 7469 26333 7481 26367
rect 7515 26333 7527 26367
rect 7469 26327 7527 26333
rect 4856 26268 5028 26296
rect 5077 26299 5135 26305
rect 4856 26256 4862 26268
rect 5077 26265 5089 26299
rect 5123 26296 5135 26299
rect 5721 26299 5779 26305
rect 5123 26268 5672 26296
rect 5123 26265 5135 26268
rect 5077 26259 5135 26265
rect 1762 26188 1768 26240
rect 1820 26188 1826 26240
rect 2774 26188 2780 26240
rect 2832 26228 2838 26240
rect 5166 26237 5172 26240
rect 2961 26231 3019 26237
rect 2961 26228 2973 26231
rect 2832 26200 2973 26228
rect 2832 26188 2838 26200
rect 2961 26197 2973 26200
rect 3007 26197 3019 26231
rect 2961 26191 3019 26197
rect 5162 26191 5172 26237
rect 5166 26188 5172 26191
rect 5224 26188 5230 26240
rect 5644 26228 5672 26268
rect 5721 26265 5733 26299
rect 5767 26296 5779 26299
rect 6270 26296 6276 26308
rect 5767 26268 6276 26296
rect 5767 26265 5779 26268
rect 5721 26259 5779 26265
rect 6270 26256 6276 26268
rect 6328 26256 6334 26308
rect 6840 26296 6868 26327
rect 6380 26268 6868 26296
rect 7116 26296 7144 26327
rect 7576 26296 7604 26540
rect 9858 26528 9864 26540
rect 9916 26528 9922 26580
rect 9950 26528 9956 26580
rect 10008 26568 10014 26580
rect 10689 26571 10747 26577
rect 10689 26568 10701 26571
rect 10008 26540 10701 26568
rect 10008 26528 10014 26540
rect 10689 26537 10701 26540
rect 10735 26537 10747 26571
rect 10689 26531 10747 26537
rect 11057 26571 11115 26577
rect 11057 26537 11069 26571
rect 11103 26568 11115 26571
rect 11146 26568 11152 26580
rect 11103 26540 11152 26568
rect 11103 26537 11115 26540
rect 11057 26531 11115 26537
rect 11146 26528 11152 26540
rect 11204 26528 11210 26580
rect 12250 26528 12256 26580
rect 12308 26568 12314 26580
rect 12526 26568 12532 26580
rect 12308 26540 12532 26568
rect 12308 26528 12314 26540
rect 12526 26528 12532 26540
rect 12584 26528 12590 26580
rect 18322 26528 18328 26580
rect 18380 26568 18386 26580
rect 19429 26571 19487 26577
rect 19429 26568 19441 26571
rect 18380 26540 19441 26568
rect 18380 26528 18386 26540
rect 19429 26537 19441 26540
rect 19475 26537 19487 26571
rect 19429 26531 19487 26537
rect 19613 26571 19671 26577
rect 19613 26537 19625 26571
rect 19659 26568 19671 26571
rect 20162 26568 20168 26580
rect 19659 26540 20168 26568
rect 19659 26537 19671 26540
rect 19613 26531 19671 26537
rect 20162 26528 20168 26540
rect 20220 26528 20226 26580
rect 22646 26528 22652 26580
rect 22704 26568 22710 26580
rect 22833 26571 22891 26577
rect 22833 26568 22845 26571
rect 22704 26540 22845 26568
rect 22704 26528 22710 26540
rect 22833 26537 22845 26540
rect 22879 26537 22891 26571
rect 22833 26531 22891 26537
rect 8496 26472 9076 26500
rect 7650 26324 7656 26376
rect 7708 26364 7714 26376
rect 8496 26373 8524 26472
rect 8588 26404 8984 26432
rect 8588 26376 8616 26404
rect 8481 26367 8539 26373
rect 8481 26364 8493 26367
rect 7708 26336 8493 26364
rect 7708 26324 7714 26336
rect 8481 26333 8493 26336
rect 8527 26333 8539 26367
rect 8481 26327 8539 26333
rect 8570 26324 8576 26376
rect 8628 26324 8634 26376
rect 8754 26324 8760 26376
rect 8812 26324 8818 26376
rect 8956 26373 8984 26404
rect 9048 26373 9076 26472
rect 10226 26460 10232 26512
rect 10284 26500 10290 26512
rect 10284 26472 10640 26500
rect 10284 26460 10290 26472
rect 9784 26404 10364 26432
rect 9784 26376 9812 26404
rect 8941 26367 8999 26373
rect 8941 26333 8953 26367
rect 8987 26333 8999 26367
rect 8941 26327 8999 26333
rect 9033 26367 9091 26373
rect 9033 26333 9045 26367
rect 9079 26333 9091 26367
rect 9033 26327 9091 26333
rect 9217 26367 9275 26373
rect 9217 26333 9229 26367
rect 9263 26333 9275 26367
rect 9217 26327 9275 26333
rect 7116 26268 7604 26296
rect 8772 26296 8800 26324
rect 9232 26296 9260 26327
rect 9766 26324 9772 26376
rect 9824 26324 9830 26376
rect 10045 26367 10103 26373
rect 10045 26333 10057 26367
rect 10091 26364 10103 26367
rect 10226 26364 10232 26376
rect 10091 26336 10232 26364
rect 10091 26333 10103 26336
rect 10045 26327 10103 26333
rect 10226 26324 10232 26336
rect 10284 26324 10290 26376
rect 10336 26373 10364 26404
rect 10321 26367 10379 26373
rect 10321 26333 10333 26367
rect 10367 26333 10379 26367
rect 10321 26327 10379 26333
rect 10502 26324 10508 26376
rect 10560 26324 10566 26376
rect 10612 26373 10640 26472
rect 11698 26460 11704 26512
rect 11756 26500 11762 26512
rect 11756 26472 13492 26500
rect 11756 26460 11762 26472
rect 11882 26392 11888 26444
rect 11940 26432 11946 26444
rect 11940 26404 13308 26432
rect 11940 26392 11946 26404
rect 10597 26367 10655 26373
rect 10597 26333 10609 26367
rect 10643 26333 10655 26367
rect 10597 26327 10655 26333
rect 8772 26268 9260 26296
rect 9953 26299 10011 26305
rect 6380 26228 6408 26268
rect 9953 26265 9965 26299
rect 9999 26296 10011 26299
rect 10612 26296 10640 26327
rect 10686 26324 10692 26376
rect 10744 26364 10750 26376
rect 10873 26367 10931 26373
rect 10873 26364 10885 26367
rect 10744 26336 10885 26364
rect 10744 26324 10750 26336
rect 10873 26333 10885 26336
rect 10919 26333 10931 26367
rect 10873 26327 10931 26333
rect 11149 26367 11207 26373
rect 11149 26333 11161 26367
rect 11195 26364 11207 26367
rect 11514 26364 11520 26376
rect 11195 26336 11520 26364
rect 11195 26333 11207 26336
rect 11149 26327 11207 26333
rect 11514 26324 11520 26336
rect 11572 26364 11578 26376
rect 12158 26364 12164 26376
rect 11572 26336 12164 26364
rect 11572 26324 11578 26336
rect 12158 26324 12164 26336
rect 12216 26324 12222 26376
rect 12250 26324 12256 26376
rect 12308 26324 12314 26376
rect 12529 26367 12587 26373
rect 12529 26333 12541 26367
rect 12575 26364 12587 26367
rect 12710 26364 12716 26376
rect 12575 26336 12716 26364
rect 12575 26333 12587 26336
rect 12529 26327 12587 26333
rect 12710 26324 12716 26336
rect 12768 26324 12774 26376
rect 12802 26324 12808 26376
rect 12860 26324 12866 26376
rect 13078 26324 13084 26376
rect 13136 26324 13142 26376
rect 13280 26373 13308 26404
rect 13464 26373 13492 26472
rect 21450 26460 21456 26512
rect 21508 26500 21514 26512
rect 22848 26500 22876 26531
rect 24210 26528 24216 26580
rect 24268 26568 24274 26580
rect 24854 26568 24860 26580
rect 24268 26540 24860 26568
rect 24268 26528 24274 26540
rect 24854 26528 24860 26540
rect 24912 26568 24918 26580
rect 25041 26571 25099 26577
rect 25041 26568 25053 26571
rect 24912 26540 25053 26568
rect 24912 26528 24918 26540
rect 25041 26537 25053 26540
rect 25087 26537 25099 26571
rect 25041 26531 25099 26537
rect 26053 26571 26111 26577
rect 26053 26537 26065 26571
rect 26099 26568 26111 26571
rect 26234 26568 26240 26580
rect 26099 26540 26240 26568
rect 26099 26537 26111 26540
rect 26053 26531 26111 26537
rect 24946 26500 24952 26512
rect 21508 26472 22094 26500
rect 22848 26472 24952 26500
rect 21508 26460 21514 26472
rect 19610 26392 19616 26444
rect 19668 26432 19674 26444
rect 20073 26435 20131 26441
rect 20073 26432 20085 26435
rect 19668 26404 20085 26432
rect 19668 26392 19674 26404
rect 20073 26401 20085 26404
rect 20119 26432 20131 26435
rect 20622 26432 20628 26444
rect 20119 26404 20628 26432
rect 20119 26401 20131 26404
rect 20073 26395 20131 26401
rect 20622 26392 20628 26404
rect 20680 26392 20686 26444
rect 21468 26432 21496 26460
rect 20732 26404 21496 26432
rect 22066 26432 22094 26472
rect 24946 26460 24952 26472
rect 25004 26460 25010 26512
rect 25056 26432 25084 26531
rect 26234 26528 26240 26540
rect 26292 26528 26298 26580
rect 26697 26571 26755 26577
rect 26697 26537 26709 26571
rect 26743 26568 26755 26571
rect 26786 26568 26792 26580
rect 26743 26540 26792 26568
rect 26743 26537 26755 26540
rect 26697 26531 26755 26537
rect 26786 26528 26792 26540
rect 26844 26528 26850 26580
rect 27706 26460 27712 26512
rect 27764 26460 27770 26512
rect 25133 26435 25191 26441
rect 25133 26432 25145 26435
rect 22066 26404 24992 26432
rect 25056 26404 25145 26432
rect 13173 26367 13231 26373
rect 13173 26333 13185 26367
rect 13219 26333 13231 26367
rect 13173 26327 13231 26333
rect 13265 26367 13323 26373
rect 13265 26333 13277 26367
rect 13311 26333 13323 26367
rect 13265 26327 13323 26333
rect 13449 26367 13507 26373
rect 13449 26333 13461 26367
rect 13495 26333 13507 26367
rect 13449 26327 13507 26333
rect 9999 26268 10640 26296
rect 9999 26265 10011 26268
rect 9953 26259 10011 26265
rect 12066 26256 12072 26308
rect 12124 26256 12130 26308
rect 13188 26296 13216 26327
rect 19978 26324 19984 26376
rect 20036 26324 20042 26376
rect 20162 26324 20168 26376
rect 20220 26364 20226 26376
rect 20257 26367 20315 26373
rect 20257 26364 20269 26367
rect 20220 26336 20269 26364
rect 20220 26324 20226 26336
rect 20257 26333 20269 26336
rect 20303 26333 20315 26367
rect 20257 26327 20315 26333
rect 13004 26268 13216 26296
rect 20272 26296 20300 26327
rect 20346 26324 20352 26376
rect 20404 26364 20410 26376
rect 20441 26367 20499 26373
rect 20441 26364 20453 26367
rect 20404 26336 20453 26364
rect 20404 26324 20410 26336
rect 20441 26333 20453 26336
rect 20487 26364 20499 26367
rect 20732 26364 20760 26404
rect 20487 26336 20760 26364
rect 20487 26333 20499 26336
rect 20441 26327 20499 26333
rect 20806 26324 20812 26376
rect 20864 26364 20870 26376
rect 20901 26367 20959 26373
rect 20901 26364 20913 26367
rect 20864 26336 20913 26364
rect 20864 26324 20870 26336
rect 20901 26333 20913 26336
rect 20947 26333 20959 26367
rect 20901 26327 20959 26333
rect 20993 26367 21051 26373
rect 20993 26333 21005 26367
rect 21039 26364 21051 26367
rect 21818 26364 21824 26376
rect 21039 26336 21824 26364
rect 21039 26333 21051 26336
rect 20993 26327 21051 26333
rect 21818 26324 21824 26336
rect 21876 26324 21882 26376
rect 23109 26367 23167 26373
rect 23109 26333 23121 26367
rect 23155 26364 23167 26367
rect 24210 26364 24216 26376
rect 23155 26336 24216 26364
rect 23155 26333 23167 26336
rect 23109 26327 23167 26333
rect 24210 26324 24216 26336
rect 24268 26324 24274 26376
rect 24854 26324 24860 26376
rect 24912 26324 24918 26376
rect 24964 26364 24992 26404
rect 25133 26401 25145 26404
rect 25179 26401 25191 26435
rect 25133 26395 25191 26401
rect 25618 26435 25676 26441
rect 25618 26401 25630 26435
rect 25664 26401 25676 26435
rect 25618 26395 25676 26401
rect 25314 26364 25320 26376
rect 24964 26336 25320 26364
rect 25314 26324 25320 26336
rect 25372 26324 25378 26376
rect 25406 26324 25412 26376
rect 25464 26364 25470 26376
rect 25501 26367 25559 26373
rect 25501 26364 25513 26367
rect 25464 26336 25513 26364
rect 25464 26324 25470 26336
rect 25501 26333 25513 26336
rect 25547 26333 25559 26367
rect 25633 26364 25661 26395
rect 25774 26364 25780 26376
rect 25633 26336 25780 26364
rect 25501 26327 25559 26333
rect 25774 26324 25780 26336
rect 25832 26324 25838 26376
rect 26513 26367 26571 26373
rect 26513 26364 26525 26367
rect 26252 26336 26525 26364
rect 20622 26296 20628 26308
rect 20272 26268 20628 26296
rect 13004 26240 13032 26268
rect 20622 26256 20628 26268
rect 20680 26296 20686 26308
rect 22462 26296 22468 26308
rect 20680 26268 22468 26296
rect 20680 26256 20686 26268
rect 22462 26256 22468 26268
rect 22520 26256 22526 26308
rect 22925 26299 22983 26305
rect 22925 26265 22937 26299
rect 22971 26296 22983 26299
rect 23014 26296 23020 26308
rect 22971 26268 23020 26296
rect 22971 26265 22983 26268
rect 22925 26259 22983 26265
rect 23014 26256 23020 26268
rect 23072 26296 23078 26308
rect 23658 26296 23664 26308
rect 23072 26268 23664 26296
rect 23072 26256 23078 26268
rect 23658 26256 23664 26268
rect 23716 26256 23722 26308
rect 24670 26256 24676 26308
rect 24728 26296 24734 26308
rect 25424 26296 25452 26324
rect 26252 26308 26280 26336
rect 26513 26333 26525 26336
rect 26559 26333 26571 26367
rect 26513 26327 26571 26333
rect 26694 26324 26700 26376
rect 26752 26324 26758 26376
rect 27522 26324 27528 26376
rect 27580 26324 27586 26376
rect 24728 26268 25452 26296
rect 26145 26299 26203 26305
rect 24728 26256 24734 26268
rect 26145 26265 26157 26299
rect 26191 26296 26203 26299
rect 26234 26296 26240 26308
rect 26191 26268 26240 26296
rect 26191 26265 26203 26268
rect 26145 26259 26203 26265
rect 26234 26256 26240 26268
rect 26292 26256 26298 26308
rect 26326 26256 26332 26308
rect 26384 26256 26390 26308
rect 5644 26200 6408 26228
rect 6546 26188 6552 26240
rect 6604 26188 6610 26240
rect 7650 26188 7656 26240
rect 7708 26188 7714 26240
rect 8662 26188 8668 26240
rect 8720 26188 8726 26240
rect 9398 26188 9404 26240
rect 9456 26188 9462 26240
rect 10042 26188 10048 26240
rect 10100 26188 10106 26240
rect 10137 26231 10195 26237
rect 10137 26197 10149 26231
rect 10183 26228 10195 26231
rect 10410 26228 10416 26240
rect 10183 26200 10416 26228
rect 10183 26197 10195 26200
rect 10137 26191 10195 26197
rect 10410 26188 10416 26200
rect 10468 26188 10474 26240
rect 10502 26188 10508 26240
rect 10560 26228 10566 26240
rect 12342 26228 12348 26240
rect 10560 26200 12348 26228
rect 10560 26188 10566 26200
rect 12342 26188 12348 26200
rect 12400 26228 12406 26240
rect 12437 26231 12495 26237
rect 12437 26228 12449 26231
rect 12400 26200 12449 26228
rect 12400 26188 12406 26200
rect 12437 26197 12449 26200
rect 12483 26197 12495 26231
rect 12437 26191 12495 26197
rect 12526 26188 12532 26240
rect 12584 26228 12590 26240
rect 12621 26231 12679 26237
rect 12621 26228 12633 26231
rect 12584 26200 12633 26228
rect 12584 26188 12590 26200
rect 12621 26197 12633 26200
rect 12667 26197 12679 26231
rect 12621 26191 12679 26197
rect 12986 26188 12992 26240
rect 13044 26188 13050 26240
rect 13170 26188 13176 26240
rect 13228 26188 13234 26240
rect 19613 26231 19671 26237
rect 19613 26197 19625 26231
rect 19659 26228 19671 26231
rect 20806 26228 20812 26240
rect 19659 26200 20812 26228
rect 19659 26197 19671 26200
rect 19613 26191 19671 26197
rect 20806 26188 20812 26200
rect 20864 26188 20870 26240
rect 24578 26188 24584 26240
rect 24636 26228 24642 26240
rect 25130 26228 25136 26240
rect 24636 26200 25136 26228
rect 24636 26188 24642 26200
rect 25130 26188 25136 26200
rect 25188 26228 25194 26240
rect 25409 26231 25467 26237
rect 25409 26228 25421 26231
rect 25188 26200 25421 26228
rect 25188 26188 25194 26200
rect 25409 26197 25421 26200
rect 25455 26197 25467 26231
rect 25409 26191 25467 26197
rect 25774 26188 25780 26240
rect 25832 26188 25838 26240
rect 1104 26138 28152 26160
rect 1104 26086 4874 26138
rect 4926 26086 4938 26138
rect 4990 26086 5002 26138
rect 5054 26086 5066 26138
rect 5118 26086 5130 26138
rect 5182 26086 28152 26138
rect 1104 26064 28152 26086
rect 2774 25984 2780 26036
rect 2832 25984 2838 26036
rect 8113 26027 8171 26033
rect 8113 25993 8125 26027
rect 8159 26024 8171 26027
rect 8570 26024 8576 26036
rect 8159 25996 8576 26024
rect 8159 25993 8171 25996
rect 8113 25987 8171 25993
rect 8570 25984 8576 25996
rect 8628 25984 8634 26036
rect 12710 25984 12716 26036
rect 12768 25984 12774 26036
rect 25774 25984 25780 26036
rect 25832 26024 25838 26036
rect 26437 26027 26495 26033
rect 26437 26024 26449 26027
rect 25832 25996 26449 26024
rect 25832 25984 25838 25996
rect 26437 25993 26449 25996
rect 26483 25993 26495 26027
rect 26437 25987 26495 25993
rect 26605 26027 26663 26033
rect 26605 25993 26617 26027
rect 26651 26024 26663 26027
rect 27522 26024 27528 26036
rect 26651 25996 27528 26024
rect 26651 25993 26663 25996
rect 26605 25987 26663 25993
rect 27522 25984 27528 25996
rect 27580 25984 27586 26036
rect 7650 25916 7656 25968
rect 7708 25956 7714 25968
rect 7745 25959 7803 25965
rect 7745 25956 7757 25959
rect 7708 25928 7757 25956
rect 7708 25916 7714 25928
rect 7745 25925 7757 25928
rect 7791 25925 7803 25959
rect 7745 25919 7803 25925
rect 10042 25916 10048 25968
rect 10100 25956 10106 25968
rect 10318 25956 10324 25968
rect 10100 25928 10324 25956
rect 10100 25916 10106 25928
rect 10318 25916 10324 25928
rect 10376 25956 10382 25968
rect 10376 25928 10640 25956
rect 10376 25916 10382 25928
rect 3053 25891 3111 25897
rect 3053 25857 3065 25891
rect 3099 25888 3111 25891
rect 3418 25888 3424 25900
rect 3099 25860 3424 25888
rect 3099 25857 3111 25860
rect 3053 25851 3111 25857
rect 3418 25848 3424 25860
rect 3476 25848 3482 25900
rect 7926 25848 7932 25900
rect 7984 25848 7990 25900
rect 10410 25848 10416 25900
rect 10468 25848 10474 25900
rect 10612 25897 10640 25928
rect 26234 25916 26240 25968
rect 26292 25956 26298 25968
rect 27154 25956 27160 25968
rect 26292 25928 27160 25956
rect 26292 25916 26298 25928
rect 27154 25916 27160 25928
rect 27212 25916 27218 25968
rect 10597 25891 10655 25897
rect 10597 25857 10609 25891
rect 10643 25857 10655 25891
rect 10597 25851 10655 25857
rect 12526 25848 12532 25900
rect 12584 25848 12590 25900
rect 12710 25848 12716 25900
rect 12768 25888 12774 25900
rect 13170 25888 13176 25900
rect 12768 25860 13176 25888
rect 12768 25848 12774 25860
rect 13170 25848 13176 25860
rect 13228 25848 13234 25900
rect 21818 25848 21824 25900
rect 21876 25888 21882 25900
rect 25774 25888 25780 25900
rect 21876 25860 25780 25888
rect 21876 25848 21882 25860
rect 25774 25848 25780 25860
rect 25832 25848 25838 25900
rect 26326 25848 26332 25900
rect 26384 25888 26390 25900
rect 26973 25891 27031 25897
rect 26973 25888 26985 25891
rect 26384 25860 26985 25888
rect 26384 25848 26390 25860
rect 26973 25857 26985 25860
rect 27019 25857 27031 25891
rect 26973 25851 27031 25857
rect 23750 25712 23756 25764
rect 23808 25752 23814 25764
rect 26970 25752 26976 25764
rect 23808 25724 26976 25752
rect 23808 25712 23814 25724
rect 26970 25712 26976 25724
rect 27028 25712 27034 25764
rect 10502 25644 10508 25696
rect 10560 25644 10566 25696
rect 20070 25644 20076 25696
rect 20128 25684 20134 25696
rect 20438 25684 20444 25696
rect 20128 25656 20444 25684
rect 20128 25644 20134 25656
rect 20438 25644 20444 25656
rect 20496 25684 20502 25696
rect 25498 25684 25504 25696
rect 20496 25656 25504 25684
rect 20496 25644 20502 25656
rect 25498 25644 25504 25656
rect 25556 25684 25562 25696
rect 25866 25684 25872 25696
rect 25556 25656 25872 25684
rect 25556 25644 25562 25656
rect 25866 25644 25872 25656
rect 25924 25644 25930 25696
rect 26418 25644 26424 25696
rect 26476 25684 26482 25696
rect 26694 25684 26700 25696
rect 26476 25656 26700 25684
rect 26476 25644 26482 25656
rect 26694 25644 26700 25656
rect 26752 25684 26758 25696
rect 27065 25687 27123 25693
rect 27065 25684 27077 25687
rect 26752 25656 27077 25684
rect 26752 25644 26758 25656
rect 27065 25653 27077 25656
rect 27111 25653 27123 25687
rect 27065 25647 27123 25653
rect 1104 25594 28152 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 28152 25594
rect 1104 25520 28152 25542
rect 20438 25440 20444 25492
rect 20496 25440 20502 25492
rect 20622 25440 20628 25492
rect 20680 25440 20686 25492
rect 20990 25440 20996 25492
rect 21048 25440 21054 25492
rect 23014 25480 23020 25492
rect 22480 25452 23020 25480
rect 7193 25415 7251 25421
rect 7193 25412 7205 25415
rect 6472 25384 7205 25412
rect 2498 25304 2504 25356
rect 2556 25304 2562 25356
rect 2774 25236 2780 25288
rect 2832 25236 2838 25288
rect 5718 25236 5724 25288
rect 5776 25276 5782 25288
rect 6472 25285 6500 25384
rect 7193 25381 7205 25384
rect 7239 25381 7251 25415
rect 7193 25375 7251 25381
rect 10042 25372 10048 25424
rect 10100 25412 10106 25424
rect 10502 25412 10508 25424
rect 10100 25384 10508 25412
rect 10100 25372 10106 25384
rect 10502 25372 10508 25384
rect 10560 25412 10566 25424
rect 10560 25384 15148 25412
rect 10560 25372 10566 25384
rect 6546 25304 6552 25356
rect 6604 25344 6610 25356
rect 6917 25347 6975 25353
rect 6917 25344 6929 25347
rect 6604 25316 6929 25344
rect 6604 25304 6610 25316
rect 6917 25313 6929 25316
rect 6963 25313 6975 25347
rect 6917 25307 6975 25313
rect 7653 25347 7711 25353
rect 7653 25313 7665 25347
rect 7699 25344 7711 25347
rect 13078 25344 13084 25356
rect 7699 25316 8064 25344
rect 7699 25313 7711 25316
rect 7653 25307 7711 25313
rect 6457 25279 6515 25285
rect 6457 25276 6469 25279
rect 5776 25248 6469 25276
rect 5776 25236 5782 25248
rect 6457 25245 6469 25248
rect 6503 25245 6515 25279
rect 6457 25239 6515 25245
rect 7558 25236 7564 25288
rect 7616 25236 7622 25288
rect 7745 25279 7803 25285
rect 7745 25245 7757 25279
rect 7791 25276 7803 25279
rect 7926 25276 7932 25288
rect 7791 25248 7932 25276
rect 7791 25245 7803 25248
rect 7745 25239 7803 25245
rect 5350 25168 5356 25220
rect 5408 25208 5414 25220
rect 7760 25208 7788 25239
rect 7926 25236 7932 25248
rect 7984 25236 7990 25288
rect 8036 25285 8064 25316
rect 12636 25316 13084 25344
rect 8021 25279 8079 25285
rect 8021 25245 8033 25279
rect 8067 25245 8079 25279
rect 8021 25239 8079 25245
rect 8205 25279 8263 25285
rect 8205 25245 8217 25279
rect 8251 25276 8263 25279
rect 8570 25276 8576 25288
rect 8251 25248 8576 25276
rect 8251 25245 8263 25248
rect 8205 25239 8263 25245
rect 8570 25236 8576 25248
rect 8628 25236 8634 25288
rect 8662 25236 8668 25288
rect 8720 25276 8726 25288
rect 9309 25279 9367 25285
rect 9309 25276 9321 25279
rect 8720 25248 9321 25276
rect 8720 25236 8726 25248
rect 9309 25245 9321 25248
rect 9355 25245 9367 25279
rect 9309 25239 9367 25245
rect 9398 25236 9404 25288
rect 9456 25276 9462 25288
rect 9493 25279 9551 25285
rect 9493 25276 9505 25279
rect 9456 25248 9505 25276
rect 9456 25236 9462 25248
rect 9493 25245 9505 25248
rect 9539 25276 9551 25279
rect 10045 25279 10103 25285
rect 10045 25276 10057 25279
rect 9539 25248 10057 25276
rect 9539 25245 9551 25248
rect 9493 25239 9551 25245
rect 10045 25245 10057 25248
rect 10091 25245 10103 25279
rect 10045 25239 10103 25245
rect 10199 25279 10257 25285
rect 10199 25245 10211 25279
rect 10245 25276 10257 25279
rect 10410 25276 10416 25288
rect 10245 25248 10416 25276
rect 10245 25245 10257 25248
rect 10199 25239 10257 25245
rect 5408 25180 7788 25208
rect 10060 25208 10088 25239
rect 10410 25236 10416 25248
rect 10468 25236 10474 25288
rect 11974 25236 11980 25288
rect 12032 25276 12038 25288
rect 12342 25276 12348 25288
rect 12032 25248 12348 25276
rect 12032 25236 12038 25248
rect 12342 25236 12348 25248
rect 12400 25236 12406 25288
rect 12434 25236 12440 25288
rect 12492 25236 12498 25288
rect 12636 25285 12664 25316
rect 13078 25304 13084 25316
rect 13136 25304 13142 25356
rect 15120 25353 15148 25384
rect 15562 25372 15568 25424
rect 15620 25412 15626 25424
rect 15620 25384 16068 25412
rect 15620 25372 15626 25384
rect 15105 25347 15163 25353
rect 15105 25313 15117 25347
rect 15151 25344 15163 25347
rect 15286 25344 15292 25356
rect 15151 25316 15292 25344
rect 15151 25313 15163 25316
rect 15105 25307 15163 25313
rect 15286 25304 15292 25316
rect 15344 25344 15350 25356
rect 15344 25316 15700 25344
rect 15344 25304 15350 25316
rect 12621 25279 12679 25285
rect 12621 25245 12633 25279
rect 12667 25245 12679 25279
rect 12621 25239 12679 25245
rect 12710 25236 12716 25288
rect 12768 25236 12774 25288
rect 15473 25279 15531 25285
rect 15473 25245 15485 25279
rect 15519 25245 15531 25279
rect 15473 25239 15531 25245
rect 15194 25208 15200 25220
rect 10060 25180 15200 25208
rect 5408 25168 5414 25180
rect 15194 25168 15200 25180
rect 15252 25208 15258 25220
rect 15488 25208 15516 25239
rect 15562 25236 15568 25288
rect 15620 25236 15626 25288
rect 15672 25276 15700 25316
rect 16040 25285 16068 25384
rect 22370 25344 22376 25356
rect 21100 25316 22376 25344
rect 15933 25279 15991 25285
rect 15672 25270 15884 25276
rect 15933 25270 15945 25279
rect 15672 25248 15945 25270
rect 15856 25245 15945 25248
rect 15979 25245 15991 25279
rect 15856 25242 15991 25245
rect 15933 25239 15991 25242
rect 16025 25279 16083 25285
rect 16025 25245 16037 25279
rect 16071 25245 16083 25279
rect 16025 25239 16083 25245
rect 16114 25236 16120 25288
rect 16172 25236 16178 25288
rect 21100 25285 21128 25316
rect 22370 25304 22376 25316
rect 22428 25304 22434 25356
rect 21085 25279 21143 25285
rect 21085 25245 21097 25279
rect 21131 25245 21143 25279
rect 21085 25239 21143 25245
rect 21818 25236 21824 25288
rect 21876 25276 21882 25288
rect 22480 25285 22508 25452
rect 23014 25440 23020 25452
rect 23072 25480 23078 25492
rect 23385 25483 23443 25489
rect 23385 25480 23397 25483
rect 23072 25452 23397 25480
rect 23072 25440 23078 25452
rect 23385 25449 23397 25452
rect 23431 25449 23443 25483
rect 23385 25443 23443 25449
rect 27154 25440 27160 25492
rect 27212 25440 27218 25492
rect 22738 25372 22744 25424
rect 22796 25412 22802 25424
rect 22925 25415 22983 25421
rect 22925 25412 22937 25415
rect 22796 25384 22937 25412
rect 22796 25372 22802 25384
rect 22925 25381 22937 25384
rect 22971 25381 22983 25415
rect 22925 25375 22983 25381
rect 24946 25372 24952 25424
rect 25004 25412 25010 25424
rect 26329 25415 26387 25421
rect 26329 25412 26341 25415
rect 25004 25384 26341 25412
rect 25004 25372 25010 25384
rect 26329 25381 26341 25384
rect 26375 25381 26387 25415
rect 26329 25375 26387 25381
rect 23290 25344 23296 25356
rect 22664 25316 23296 25344
rect 22664 25288 22692 25316
rect 23290 25304 23296 25316
rect 23348 25304 23354 25356
rect 25958 25344 25964 25356
rect 25792 25316 25964 25344
rect 22465 25279 22523 25285
rect 22465 25276 22477 25279
rect 21876 25248 22477 25276
rect 21876 25236 21882 25248
rect 22465 25245 22477 25248
rect 22511 25245 22523 25279
rect 22465 25239 22523 25245
rect 22646 25236 22652 25288
rect 22704 25236 22710 25288
rect 22833 25279 22891 25285
rect 22833 25245 22845 25279
rect 22879 25276 22891 25279
rect 23201 25279 23259 25285
rect 23201 25276 23213 25279
rect 22879 25248 23213 25276
rect 22879 25245 22891 25248
rect 22833 25239 22891 25245
rect 23201 25245 23213 25248
rect 23247 25276 23259 25279
rect 23382 25276 23388 25288
rect 23247 25248 23388 25276
rect 23247 25245 23259 25248
rect 23201 25239 23259 25245
rect 23382 25236 23388 25248
rect 23440 25236 23446 25288
rect 25792 25285 25820 25316
rect 25958 25304 25964 25316
rect 26016 25304 26022 25356
rect 26145 25347 26203 25353
rect 26145 25313 26157 25347
rect 26191 25344 26203 25347
rect 26191 25316 27568 25344
rect 26191 25313 26203 25316
rect 26145 25307 26203 25313
rect 25777 25279 25835 25285
rect 25777 25245 25789 25279
rect 25823 25245 25835 25279
rect 25777 25239 25835 25245
rect 25866 25236 25872 25288
rect 25924 25236 25930 25288
rect 26234 25236 26240 25288
rect 26292 25236 26298 25288
rect 27540 25285 27568 25316
rect 26513 25279 26571 25285
rect 26513 25245 26525 25279
rect 26559 25245 26571 25279
rect 26513 25239 26571 25245
rect 27525 25279 27583 25285
rect 27525 25245 27537 25279
rect 27571 25245 27583 25279
rect 27525 25239 27583 25245
rect 15252 25180 15516 25208
rect 15749 25211 15807 25217
rect 15252 25168 15258 25180
rect 15749 25177 15761 25211
rect 15795 25208 15807 25211
rect 16666 25208 16672 25220
rect 15795 25180 16672 25208
rect 15795 25177 15807 25180
rect 15749 25171 15807 25177
rect 16666 25168 16672 25180
rect 16724 25168 16730 25220
rect 20806 25168 20812 25220
rect 20864 25168 20870 25220
rect 22186 25168 22192 25220
rect 22244 25208 22250 25220
rect 22925 25211 22983 25217
rect 22925 25208 22937 25211
rect 22244 25180 22937 25208
rect 22244 25168 22250 25180
rect 22925 25177 22937 25180
rect 22971 25208 22983 25211
rect 23014 25208 23020 25220
rect 22971 25180 23020 25208
rect 22971 25177 22983 25180
rect 22925 25171 22983 25177
rect 23014 25168 23020 25180
rect 23072 25168 23078 25220
rect 23109 25211 23167 25217
rect 23109 25177 23121 25211
rect 23155 25208 23167 25211
rect 23477 25211 23535 25217
rect 23155 25180 23428 25208
rect 23155 25177 23167 25180
rect 23109 25171 23167 25177
rect 3421 25143 3479 25149
rect 3421 25109 3433 25143
rect 3467 25140 3479 25143
rect 3510 25140 3516 25152
rect 3467 25112 3516 25140
rect 3467 25109 3479 25112
rect 3421 25103 3479 25109
rect 3510 25100 3516 25112
rect 3568 25100 3574 25152
rect 6825 25143 6883 25149
rect 6825 25109 6837 25143
rect 6871 25140 6883 25143
rect 7282 25140 7288 25152
rect 6871 25112 7288 25140
rect 6871 25109 6883 25112
rect 6825 25103 6883 25109
rect 7282 25100 7288 25112
rect 7340 25100 7346 25152
rect 7374 25100 7380 25152
rect 7432 25100 7438 25152
rect 8205 25143 8263 25149
rect 8205 25109 8217 25143
rect 8251 25140 8263 25143
rect 8386 25140 8392 25152
rect 8251 25112 8392 25140
rect 8251 25109 8263 25112
rect 8205 25103 8263 25109
rect 8386 25100 8392 25112
rect 8444 25100 8450 25152
rect 9490 25100 9496 25152
rect 9548 25100 9554 25152
rect 10413 25143 10471 25149
rect 10413 25109 10425 25143
rect 10459 25140 10471 25143
rect 10502 25140 10508 25152
rect 10459 25112 10508 25140
rect 10459 25109 10471 25112
rect 10413 25103 10471 25109
rect 10502 25100 10508 25112
rect 10560 25100 10566 25152
rect 12894 25100 12900 25152
rect 12952 25100 12958 25152
rect 16301 25143 16359 25149
rect 16301 25109 16313 25143
rect 16347 25140 16359 25143
rect 16758 25140 16764 25152
rect 16347 25112 16764 25140
rect 16347 25109 16359 25112
rect 16301 25103 16359 25109
rect 16758 25100 16764 25112
rect 16816 25100 16822 25152
rect 20609 25143 20667 25149
rect 20609 25109 20621 25143
rect 20655 25140 20667 25143
rect 20990 25140 20996 25152
rect 20655 25112 20996 25140
rect 20655 25109 20667 25112
rect 20609 25103 20667 25109
rect 20990 25100 20996 25112
rect 21048 25100 21054 25152
rect 23400 25140 23428 25180
rect 23477 25177 23489 25211
rect 23523 25208 23535 25211
rect 23566 25208 23572 25220
rect 23523 25180 23572 25208
rect 23523 25177 23535 25180
rect 23477 25171 23535 25177
rect 23566 25168 23572 25180
rect 23624 25168 23630 25220
rect 24762 25168 24768 25220
rect 24820 25208 24826 25220
rect 25593 25211 25651 25217
rect 25593 25208 25605 25211
rect 24820 25180 25605 25208
rect 24820 25168 24826 25180
rect 25593 25177 25605 25180
rect 25639 25208 25651 25211
rect 25961 25211 26019 25217
rect 25639 25180 25912 25208
rect 25639 25177 25651 25180
rect 25593 25171 25651 25177
rect 23658 25140 23664 25152
rect 23400 25112 23664 25140
rect 23658 25100 23664 25112
rect 23716 25100 23722 25152
rect 25884 25140 25912 25180
rect 25961 25177 25973 25211
rect 26007 25208 26019 25211
rect 26418 25208 26424 25220
rect 26007 25180 26424 25208
rect 26007 25177 26019 25180
rect 25961 25171 26019 25177
rect 26418 25168 26424 25180
rect 26476 25168 26482 25220
rect 26528 25152 26556 25239
rect 26697 25211 26755 25217
rect 26697 25177 26709 25211
rect 26743 25208 26755 25211
rect 26789 25211 26847 25217
rect 26789 25208 26801 25211
rect 26743 25180 26801 25208
rect 26743 25177 26755 25180
rect 26697 25171 26755 25177
rect 26789 25177 26801 25180
rect 26835 25177 26847 25211
rect 26789 25171 26847 25177
rect 26973 25211 27031 25217
rect 26973 25177 26985 25211
rect 27019 25208 27031 25211
rect 27154 25208 27160 25220
rect 27019 25180 27160 25208
rect 27019 25177 27031 25180
rect 26973 25171 27031 25177
rect 27154 25168 27160 25180
rect 27212 25168 27218 25220
rect 26510 25140 26516 25152
rect 25884 25112 26516 25140
rect 26510 25100 26516 25112
rect 26568 25100 26574 25152
rect 27706 25100 27712 25152
rect 27764 25100 27770 25152
rect 1104 25050 28152 25072
rect 1104 24998 4874 25050
rect 4926 24998 4938 25050
rect 4990 24998 5002 25050
rect 5054 24998 5066 25050
rect 5118 24998 5130 25050
rect 5182 24998 28152 25050
rect 1104 24976 28152 24998
rect 11974 24896 11980 24948
rect 12032 24936 12038 24948
rect 12069 24939 12127 24945
rect 12069 24936 12081 24939
rect 12032 24908 12081 24936
rect 12032 24896 12038 24908
rect 12069 24905 12081 24908
rect 12115 24905 12127 24939
rect 12069 24899 12127 24905
rect 12158 24896 12164 24948
rect 12216 24896 12222 24948
rect 16666 24896 16672 24948
rect 16724 24936 16730 24948
rect 17421 24939 17479 24945
rect 17421 24936 17433 24939
rect 16724 24908 17433 24936
rect 16724 24896 16730 24908
rect 17421 24905 17433 24908
rect 17467 24905 17479 24939
rect 17421 24899 17479 24905
rect 20732 24908 22968 24936
rect 10042 24828 10048 24880
rect 10100 24828 10106 24880
rect 12176 24868 12204 24896
rect 12897 24871 12955 24877
rect 12176 24840 12296 24868
rect 4249 24803 4307 24809
rect 4249 24769 4261 24803
rect 4295 24800 4307 24803
rect 5350 24800 5356 24812
rect 4295 24772 5356 24800
rect 4295 24769 4307 24772
rect 4249 24763 4307 24769
rect 5350 24760 5356 24772
rect 5408 24760 5414 24812
rect 7374 24760 7380 24812
rect 7432 24800 7438 24812
rect 7929 24803 7987 24809
rect 7929 24800 7941 24803
rect 7432 24772 7941 24800
rect 7432 24760 7438 24772
rect 7929 24769 7941 24772
rect 7975 24769 7987 24803
rect 7929 24763 7987 24769
rect 3602 24692 3608 24744
rect 3660 24732 3666 24744
rect 4157 24735 4215 24741
rect 4157 24732 4169 24735
rect 3660 24704 4169 24732
rect 3660 24692 3666 24704
rect 4157 24701 4169 24704
rect 4203 24701 4215 24735
rect 4157 24695 4215 24701
rect 4341 24735 4399 24741
rect 4341 24701 4353 24735
rect 4387 24701 4399 24735
rect 4341 24695 4399 24701
rect 4433 24735 4491 24741
rect 4433 24701 4445 24735
rect 4479 24732 4491 24735
rect 4614 24732 4620 24744
rect 4479 24704 4620 24732
rect 4479 24701 4491 24704
rect 4433 24695 4491 24701
rect 4356 24664 4384 24695
rect 4614 24692 4620 24704
rect 4672 24692 4678 24744
rect 7944 24732 7972 24763
rect 8110 24760 8116 24812
rect 8168 24760 8174 24812
rect 8386 24760 8392 24812
rect 8444 24800 8450 24812
rect 8757 24803 8815 24809
rect 8757 24800 8769 24803
rect 8444 24772 8769 24800
rect 8444 24760 8450 24772
rect 8757 24769 8769 24772
rect 8803 24769 8815 24803
rect 8757 24763 8815 24769
rect 9490 24760 9496 24812
rect 9548 24800 9554 24812
rect 9861 24803 9919 24809
rect 9861 24800 9873 24803
rect 9548 24772 9873 24800
rect 9548 24760 9554 24772
rect 9861 24769 9873 24772
rect 9907 24769 9919 24803
rect 9861 24763 9919 24769
rect 10318 24760 10324 24812
rect 10376 24760 10382 24812
rect 10502 24760 10508 24812
rect 10560 24760 10566 24812
rect 10597 24803 10655 24809
rect 10597 24769 10609 24803
rect 10643 24769 10655 24803
rect 10597 24763 10655 24769
rect 10689 24803 10747 24809
rect 10689 24769 10701 24803
rect 10735 24769 10747 24803
rect 10689 24763 10747 24769
rect 8849 24735 8907 24741
rect 8849 24732 8861 24735
rect 7944 24704 8861 24732
rect 8849 24701 8861 24704
rect 8895 24701 8907 24735
rect 8849 24695 8907 24701
rect 8941 24735 8999 24741
rect 8941 24701 8953 24735
rect 8987 24701 8999 24735
rect 8941 24695 8999 24701
rect 4798 24664 4804 24676
rect 4356 24636 4804 24664
rect 4798 24624 4804 24636
rect 4856 24624 4862 24676
rect 8110 24624 8116 24676
rect 8168 24664 8174 24676
rect 8956 24664 8984 24695
rect 10410 24692 10416 24744
rect 10468 24732 10474 24744
rect 10612 24732 10640 24763
rect 10468 24704 10640 24732
rect 10468 24692 10474 24704
rect 10704 24664 10732 24763
rect 11790 24760 11796 24812
rect 11848 24760 11854 24812
rect 12066 24760 12072 24812
rect 12124 24800 12130 24812
rect 12268 24809 12296 24840
rect 12897 24837 12909 24871
rect 12943 24868 12955 24871
rect 13078 24868 13084 24880
rect 12943 24840 13084 24868
rect 12943 24837 12955 24840
rect 12897 24831 12955 24837
rect 12161 24803 12219 24809
rect 12161 24800 12173 24803
rect 12124 24772 12173 24800
rect 12124 24760 12130 24772
rect 12161 24769 12173 24772
rect 12207 24769 12219 24803
rect 12161 24763 12219 24769
rect 12253 24803 12311 24809
rect 12253 24769 12265 24803
rect 12299 24769 12311 24803
rect 12713 24803 12771 24809
rect 12713 24800 12725 24803
rect 12253 24763 12311 24769
rect 12406 24772 12725 24800
rect 10965 24735 11023 24741
rect 10965 24701 10977 24735
rect 11011 24732 11023 24735
rect 11609 24735 11667 24741
rect 11609 24732 11621 24735
rect 11011 24704 11621 24732
rect 11011 24701 11023 24704
rect 10965 24695 11023 24701
rect 11609 24701 11621 24704
rect 11655 24732 11667 24735
rect 11974 24732 11980 24744
rect 11655 24704 11980 24732
rect 11655 24701 11667 24704
rect 11609 24695 11667 24701
rect 11974 24692 11980 24704
rect 12032 24692 12038 24744
rect 12406 24732 12434 24772
rect 12713 24769 12725 24772
rect 12759 24769 12771 24803
rect 12713 24763 12771 24769
rect 12084 24704 12434 24732
rect 12529 24735 12587 24741
rect 8168 24636 8984 24664
rect 10244 24636 10732 24664
rect 8168 24624 8174 24636
rect 4617 24599 4675 24605
rect 4617 24565 4629 24599
rect 4663 24596 4675 24599
rect 5166 24596 5172 24608
rect 4663 24568 5172 24596
rect 4663 24565 4675 24568
rect 4617 24559 4675 24565
rect 5166 24556 5172 24568
rect 5224 24556 5230 24608
rect 8570 24556 8576 24608
rect 8628 24556 8634 24608
rect 9125 24599 9183 24605
rect 9125 24565 9137 24599
rect 9171 24596 9183 24599
rect 9398 24596 9404 24608
rect 9171 24568 9404 24596
rect 9171 24565 9183 24568
rect 9125 24559 9183 24565
rect 9398 24556 9404 24568
rect 9456 24556 9462 24608
rect 9950 24556 9956 24608
rect 10008 24596 10014 24608
rect 10244 24605 10272 24636
rect 10229 24599 10287 24605
rect 10229 24596 10241 24599
rect 10008 24568 10241 24596
rect 10008 24556 10014 24568
rect 10229 24565 10241 24568
rect 10275 24565 10287 24599
rect 10229 24559 10287 24565
rect 10318 24556 10324 24608
rect 10376 24596 10382 24608
rect 12084 24596 12112 24704
rect 12529 24701 12541 24735
rect 12575 24732 12587 24735
rect 12912 24732 12940 24831
rect 13078 24828 13084 24840
rect 13136 24868 13142 24880
rect 13354 24868 13360 24880
rect 13136 24840 13360 24868
rect 13136 24828 13142 24840
rect 13354 24828 13360 24840
rect 13412 24828 13418 24880
rect 17221 24871 17279 24877
rect 17221 24868 17233 24871
rect 15304 24840 15884 24868
rect 15304 24812 15332 24840
rect 12989 24803 13047 24809
rect 12989 24769 13001 24803
rect 13035 24769 13047 24803
rect 12989 24763 13047 24769
rect 12575 24704 12940 24732
rect 12575 24701 12587 24704
rect 12529 24695 12587 24701
rect 12342 24624 12348 24676
rect 12400 24664 12406 24676
rect 13004 24664 13032 24763
rect 13170 24760 13176 24812
rect 13228 24760 13234 24812
rect 14090 24760 14096 24812
rect 14148 24800 14154 24812
rect 15013 24803 15071 24809
rect 15013 24800 15025 24803
rect 14148 24772 15025 24800
rect 14148 24760 14154 24772
rect 15013 24769 15025 24772
rect 15059 24769 15071 24803
rect 15013 24763 15071 24769
rect 15105 24803 15163 24809
rect 15105 24769 15117 24803
rect 15151 24800 15163 24803
rect 15194 24800 15200 24812
rect 15151 24772 15200 24800
rect 15151 24769 15163 24772
rect 15105 24763 15163 24769
rect 12400 24636 13032 24664
rect 15028 24664 15056 24763
rect 15194 24760 15200 24772
rect 15252 24760 15258 24812
rect 15286 24760 15292 24812
rect 15344 24760 15350 24812
rect 15562 24760 15568 24812
rect 15620 24760 15626 24812
rect 15856 24809 15884 24840
rect 16592 24840 17233 24868
rect 16592 24812 16620 24840
rect 15749 24803 15807 24809
rect 15749 24769 15761 24803
rect 15795 24769 15807 24803
rect 15749 24763 15807 24769
rect 15841 24803 15899 24809
rect 15841 24769 15853 24803
rect 15887 24769 15899 24803
rect 15841 24763 15899 24769
rect 15212 24732 15240 24760
rect 15764 24732 15792 24763
rect 16298 24760 16304 24812
rect 16356 24760 16362 24812
rect 16485 24803 16543 24809
rect 16485 24769 16497 24803
rect 16531 24800 16543 24803
rect 16574 24800 16580 24812
rect 16531 24772 16580 24800
rect 16531 24769 16543 24772
rect 16485 24763 16543 24769
rect 16574 24760 16580 24772
rect 16632 24760 16638 24812
rect 16666 24760 16672 24812
rect 16724 24760 16730 24812
rect 16758 24760 16764 24812
rect 16816 24760 16822 24812
rect 16960 24809 16988 24840
rect 17221 24837 17233 24840
rect 17267 24837 17279 24871
rect 17221 24831 17279 24837
rect 16945 24803 17003 24809
rect 16945 24769 16957 24803
rect 16991 24769 17003 24803
rect 16945 24763 17003 24769
rect 20622 24760 20628 24812
rect 20680 24800 20686 24812
rect 20732 24800 20760 24908
rect 22646 24868 22652 24880
rect 22020 24840 22652 24868
rect 20680 24772 20760 24800
rect 20680 24760 20686 24772
rect 21726 24760 21732 24812
rect 21784 24800 21790 24812
rect 21913 24803 21971 24809
rect 21913 24800 21925 24803
rect 21784 24772 21925 24800
rect 21784 24760 21790 24772
rect 21913 24769 21925 24772
rect 21959 24800 21971 24803
rect 22020 24800 22048 24840
rect 22646 24828 22652 24840
rect 22704 24828 22710 24880
rect 22940 24868 22968 24908
rect 22940 24840 23046 24868
rect 24946 24828 24952 24880
rect 25004 24868 25010 24880
rect 26145 24871 26203 24877
rect 26145 24868 26157 24871
rect 25004 24840 25544 24868
rect 25004 24828 25010 24840
rect 22281 24803 22339 24809
rect 22281 24800 22293 24803
rect 21959 24772 22048 24800
rect 22112 24772 22293 24800
rect 21959 24769 21971 24772
rect 21913 24763 21971 24769
rect 16114 24732 16120 24744
rect 15212 24704 16120 24732
rect 16114 24692 16120 24704
rect 16172 24692 16178 24744
rect 15562 24664 15568 24676
rect 15028 24636 15568 24664
rect 12400 24624 12406 24636
rect 15562 24624 15568 24636
rect 15620 24624 15626 24676
rect 16776 24664 16804 24760
rect 17129 24735 17187 24741
rect 17129 24701 17141 24735
rect 17175 24732 17187 24735
rect 17494 24732 17500 24744
rect 17175 24704 17500 24732
rect 17175 24701 17187 24704
rect 17129 24695 17187 24701
rect 17494 24692 17500 24704
rect 17552 24692 17558 24744
rect 22112 24732 22140 24772
rect 22281 24769 22293 24772
rect 22327 24769 22339 24803
rect 22281 24763 22339 24769
rect 24762 24760 24768 24812
rect 24820 24800 24826 24812
rect 25516 24809 25544 24840
rect 25976 24840 26157 24868
rect 25225 24803 25283 24809
rect 25225 24800 25237 24803
rect 24820 24772 25237 24800
rect 24820 24760 24826 24772
rect 25225 24769 25237 24772
rect 25271 24769 25283 24803
rect 25225 24763 25283 24769
rect 25501 24803 25559 24809
rect 25501 24769 25513 24803
rect 25547 24800 25559 24803
rect 25866 24800 25872 24812
rect 25547 24772 25872 24800
rect 25547 24769 25559 24772
rect 25501 24763 25559 24769
rect 25866 24760 25872 24772
rect 25924 24760 25930 24812
rect 21928 24704 22140 24732
rect 21928 24676 21956 24704
rect 22186 24692 22192 24744
rect 22244 24692 22250 24744
rect 22557 24735 22615 24741
rect 22557 24732 22569 24735
rect 22296 24704 22569 24732
rect 16776 24636 17448 24664
rect 10376 24568 12112 24596
rect 10376 24556 10382 24568
rect 12434 24556 12440 24608
rect 12492 24556 12498 24608
rect 13078 24556 13084 24608
rect 13136 24596 13142 24608
rect 13173 24599 13231 24605
rect 13173 24596 13185 24599
rect 13136 24568 13185 24596
rect 13136 24556 13142 24568
rect 13173 24565 13185 24568
rect 13219 24565 13231 24599
rect 13173 24559 13231 24565
rect 15473 24599 15531 24605
rect 15473 24565 15485 24599
rect 15519 24596 15531 24599
rect 15746 24596 15752 24608
rect 15519 24568 15752 24596
rect 15519 24565 15531 24568
rect 15473 24559 15531 24565
rect 15746 24556 15752 24568
rect 15804 24556 15810 24608
rect 15841 24599 15899 24605
rect 15841 24565 15853 24599
rect 15887 24596 15899 24599
rect 15930 24596 15936 24608
rect 15887 24568 15936 24596
rect 15887 24565 15899 24568
rect 15841 24559 15899 24565
rect 15930 24556 15936 24568
rect 15988 24556 15994 24608
rect 16393 24599 16451 24605
rect 16393 24565 16405 24599
rect 16439 24596 16451 24599
rect 17310 24596 17316 24608
rect 16439 24568 17316 24596
rect 16439 24565 16451 24568
rect 16393 24559 16451 24565
rect 17310 24556 17316 24568
rect 17368 24556 17374 24608
rect 17420 24605 17448 24636
rect 21910 24624 21916 24676
rect 21968 24624 21974 24676
rect 22002 24624 22008 24676
rect 22060 24624 22066 24676
rect 17405 24599 17463 24605
rect 17405 24565 17417 24599
rect 17451 24565 17463 24599
rect 17405 24559 17463 24565
rect 17589 24599 17647 24605
rect 17589 24565 17601 24599
rect 17635 24596 17647 24599
rect 17770 24596 17776 24608
rect 17635 24568 17776 24596
rect 17635 24565 17647 24568
rect 17589 24559 17647 24565
rect 17770 24556 17776 24568
rect 17828 24556 17834 24608
rect 22097 24599 22155 24605
rect 22097 24565 22109 24599
rect 22143 24596 22155 24599
rect 22296 24596 22324 24704
rect 22557 24701 22569 24704
rect 22603 24701 22615 24735
rect 22557 24695 22615 24701
rect 23842 24692 23848 24744
rect 23900 24732 23906 24744
rect 24029 24735 24087 24741
rect 24029 24732 24041 24735
rect 23900 24704 24041 24732
rect 23900 24692 23906 24704
rect 24029 24701 24041 24704
rect 24075 24732 24087 24735
rect 24854 24732 24860 24744
rect 24075 24704 24860 24732
rect 24075 24701 24087 24704
rect 24029 24695 24087 24701
rect 24854 24692 24860 24704
rect 24912 24692 24918 24744
rect 24946 24692 24952 24744
rect 25004 24732 25010 24744
rect 25130 24732 25136 24744
rect 25004 24704 25136 24732
rect 25004 24692 25010 24704
rect 25130 24692 25136 24704
rect 25188 24732 25194 24744
rect 25409 24735 25467 24741
rect 25409 24732 25421 24735
rect 25188 24704 25421 24732
rect 25188 24692 25194 24704
rect 25409 24701 25421 24704
rect 25455 24732 25467 24735
rect 25976 24732 26004 24840
rect 26145 24837 26157 24840
rect 26191 24868 26203 24871
rect 26786 24868 26792 24880
rect 26191 24840 26792 24868
rect 26191 24837 26203 24840
rect 26145 24831 26203 24837
rect 26786 24828 26792 24840
rect 26844 24828 26850 24880
rect 27080 24840 27292 24868
rect 26605 24803 26663 24809
rect 26605 24800 26617 24803
rect 26252 24772 26617 24800
rect 25455 24704 26004 24732
rect 25455 24701 25467 24704
rect 25409 24695 25467 24701
rect 26050 24692 26056 24744
rect 26108 24732 26114 24744
rect 26252 24732 26280 24772
rect 26605 24769 26617 24772
rect 26651 24769 26663 24803
rect 26605 24763 26663 24769
rect 26970 24760 26976 24812
rect 27028 24760 27034 24812
rect 27080 24809 27108 24840
rect 27065 24803 27123 24809
rect 27065 24769 27077 24803
rect 27111 24769 27123 24803
rect 27065 24763 27123 24769
rect 27157 24803 27215 24809
rect 27157 24769 27169 24803
rect 27203 24769 27215 24803
rect 27264 24800 27292 24840
rect 27525 24803 27583 24809
rect 27525 24800 27537 24803
rect 27264 24772 27537 24800
rect 27157 24763 27215 24769
rect 27525 24769 27537 24772
rect 27571 24769 27583 24803
rect 27525 24763 27583 24769
rect 26108 24704 26280 24732
rect 26108 24692 26114 24704
rect 26510 24692 26516 24744
rect 26568 24692 26574 24744
rect 25501 24667 25559 24673
rect 25501 24633 25513 24667
rect 25547 24664 25559 24667
rect 25777 24667 25835 24673
rect 25777 24664 25789 24667
rect 25547 24636 25789 24664
rect 25547 24633 25559 24636
rect 25501 24627 25559 24633
rect 25777 24633 25789 24636
rect 25823 24664 25835 24667
rect 26789 24667 26847 24673
rect 25823 24636 26372 24664
rect 25823 24633 25835 24636
rect 25777 24627 25835 24633
rect 22143 24568 22324 24596
rect 22143 24565 22155 24568
rect 22097 24559 22155 24565
rect 25590 24556 25596 24608
rect 25648 24556 25654 24608
rect 25866 24556 25872 24608
rect 25924 24596 25930 24608
rect 26237 24599 26295 24605
rect 26237 24596 26249 24599
rect 25924 24568 26249 24596
rect 25924 24556 25930 24568
rect 26237 24565 26249 24568
rect 26283 24565 26295 24599
rect 26344 24596 26372 24636
rect 26789 24633 26801 24667
rect 26835 24664 26847 24667
rect 27172 24664 27200 24763
rect 26835 24636 27200 24664
rect 26835 24633 26847 24636
rect 26789 24627 26847 24633
rect 27154 24596 27160 24608
rect 26344 24568 27160 24596
rect 26237 24559 26295 24565
rect 27154 24556 27160 24568
rect 27212 24556 27218 24608
rect 27706 24556 27712 24608
rect 27764 24556 27770 24608
rect 1104 24506 28152 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 28152 24506
rect 1104 24432 28152 24454
rect 3602 24352 3608 24404
rect 3660 24352 3666 24404
rect 5350 24352 5356 24404
rect 5408 24352 5414 24404
rect 7561 24395 7619 24401
rect 7561 24361 7573 24395
rect 7607 24392 7619 24395
rect 8110 24392 8116 24404
rect 7607 24364 8116 24392
rect 7607 24361 7619 24364
rect 7561 24355 7619 24361
rect 8110 24352 8116 24364
rect 8168 24352 8174 24404
rect 11974 24352 11980 24404
rect 12032 24352 12038 24404
rect 12161 24395 12219 24401
rect 12161 24361 12173 24395
rect 12207 24392 12219 24395
rect 13170 24392 13176 24404
rect 12207 24364 13176 24392
rect 12207 24361 12219 24364
rect 12161 24355 12219 24361
rect 13170 24352 13176 24364
rect 13228 24352 13234 24404
rect 16206 24352 16212 24404
rect 16264 24392 16270 24404
rect 18138 24392 18144 24404
rect 16264 24364 18144 24392
rect 16264 24352 16270 24364
rect 18138 24352 18144 24364
rect 18196 24352 18202 24404
rect 18598 24352 18604 24404
rect 18656 24392 18662 24404
rect 20993 24395 21051 24401
rect 20993 24392 21005 24395
rect 18656 24364 21005 24392
rect 18656 24352 18662 24364
rect 20993 24361 21005 24364
rect 21039 24361 21051 24395
rect 20993 24355 21051 24361
rect 21726 24352 21732 24404
rect 21784 24352 21790 24404
rect 21818 24352 21824 24404
rect 21876 24352 21882 24404
rect 22002 24352 22008 24404
rect 22060 24392 22066 24404
rect 22060 24364 23244 24392
rect 22060 24352 22066 24364
rect 4062 24324 4068 24336
rect 3068 24296 4068 24324
rect 3068 24200 3096 24296
rect 4062 24284 4068 24296
rect 4120 24284 4126 24336
rect 9306 24284 9312 24336
rect 9364 24324 9370 24336
rect 10137 24327 10195 24333
rect 10137 24324 10149 24327
rect 9364 24296 10149 24324
rect 9364 24284 9370 24296
rect 10137 24293 10149 24296
rect 10183 24293 10195 24327
rect 10137 24287 10195 24293
rect 10505 24327 10563 24333
rect 10505 24293 10517 24327
rect 10551 24324 10563 24327
rect 10551 24296 14320 24324
rect 10551 24293 10563 24296
rect 10505 24287 10563 24293
rect 3510 24216 3516 24268
rect 3568 24256 3574 24268
rect 3568 24228 4016 24256
rect 3568 24216 3574 24228
rect 842 24148 848 24200
rect 900 24188 906 24200
rect 1397 24191 1455 24197
rect 1397 24188 1409 24191
rect 900 24160 1409 24188
rect 900 24148 906 24160
rect 1397 24157 1409 24160
rect 1443 24157 1455 24191
rect 1397 24151 1455 24157
rect 1762 24148 1768 24200
rect 1820 24148 1826 24200
rect 2590 24188 2596 24200
rect 2438 24160 2596 24188
rect 2590 24148 2596 24160
rect 2648 24148 2654 24200
rect 2869 24191 2927 24197
rect 2869 24188 2881 24191
rect 2746 24160 2881 24188
rect 2498 24080 2504 24132
rect 2556 24120 2562 24132
rect 2746 24120 2774 24160
rect 2869 24157 2881 24160
rect 2915 24157 2927 24191
rect 2869 24151 2927 24157
rect 3050 24148 3056 24200
rect 3108 24148 3114 24200
rect 3620 24197 3648 24228
rect 3421 24191 3479 24197
rect 3421 24157 3433 24191
rect 3467 24157 3479 24191
rect 3421 24151 3479 24157
rect 3605 24191 3663 24197
rect 3605 24157 3617 24191
rect 3651 24157 3663 24191
rect 3605 24151 3663 24157
rect 3881 24191 3939 24197
rect 3881 24157 3893 24191
rect 3927 24157 3939 24191
rect 3988 24174 4016 24228
rect 4798 24216 4804 24268
rect 4856 24256 4862 24268
rect 7193 24259 7251 24265
rect 7193 24256 7205 24259
rect 4856 24228 7205 24256
rect 4856 24216 4862 24228
rect 7193 24225 7205 24228
rect 7239 24256 7251 24259
rect 7466 24256 7472 24268
rect 7239 24228 7472 24256
rect 7239 24225 7251 24228
rect 7193 24219 7251 24225
rect 7466 24216 7472 24228
rect 7524 24216 7530 24268
rect 9953 24259 10011 24265
rect 9692 24228 9904 24256
rect 3881 24151 3939 24157
rect 2556 24092 2774 24120
rect 2961 24123 3019 24129
rect 2556 24080 2562 24092
rect 2961 24089 2973 24123
rect 3007 24120 3019 24123
rect 3436 24120 3464 24151
rect 3896 24120 3924 24151
rect 4706 24148 4712 24200
rect 4764 24188 4770 24200
rect 4985 24191 5043 24197
rect 4985 24188 4997 24191
rect 4764 24160 4997 24188
rect 4764 24148 4770 24160
rect 4985 24157 4997 24160
rect 5031 24157 5043 24191
rect 4985 24151 5043 24157
rect 5166 24148 5172 24200
rect 5224 24148 5230 24200
rect 5261 24191 5319 24197
rect 5261 24157 5273 24191
rect 5307 24157 5319 24191
rect 5261 24151 5319 24157
rect 3007 24092 3924 24120
rect 3007 24089 3019 24092
rect 2961 24083 3019 24089
rect 4430 24080 4436 24132
rect 4488 24120 4494 24132
rect 4617 24123 4675 24129
rect 4617 24120 4629 24123
rect 4488 24092 4629 24120
rect 4488 24080 4494 24092
rect 4617 24089 4629 24092
rect 4663 24089 4675 24123
rect 4617 24083 4675 24089
rect 4890 24080 4896 24132
rect 4948 24120 4954 24132
rect 5276 24120 5304 24151
rect 7282 24148 7288 24200
rect 7340 24188 7346 24200
rect 7377 24191 7435 24197
rect 7377 24188 7389 24191
rect 7340 24160 7389 24188
rect 7340 24148 7346 24160
rect 7377 24157 7389 24160
rect 7423 24157 7435 24191
rect 7377 24151 7435 24157
rect 8570 24148 8576 24200
rect 8628 24188 8634 24200
rect 9398 24197 9404 24200
rect 9125 24191 9183 24197
rect 9125 24188 9137 24191
rect 8628 24160 9137 24188
rect 8628 24148 8634 24160
rect 9125 24157 9137 24160
rect 9171 24157 9183 24191
rect 9391 24191 9404 24197
rect 9391 24188 9403 24191
rect 9125 24151 9183 24157
rect 9324 24160 9403 24188
rect 4948 24092 5304 24120
rect 8941 24123 8999 24129
rect 4948 24080 4954 24092
rect 8941 24089 8953 24123
rect 8987 24120 8999 24123
rect 9324 24120 9352 24160
rect 9391 24157 9403 24160
rect 9391 24151 9404 24157
rect 9398 24148 9404 24151
rect 9456 24148 9462 24200
rect 9490 24148 9496 24200
rect 9548 24148 9554 24200
rect 9692 24197 9720 24228
rect 9876 24200 9904 24228
rect 9953 24225 9965 24259
rect 9999 24256 10011 24259
rect 13725 24259 13783 24265
rect 9999 24228 12204 24256
rect 9999 24225 10011 24228
rect 9953 24219 10011 24225
rect 9677 24191 9735 24197
rect 9677 24157 9689 24191
rect 9723 24157 9735 24191
rect 9677 24151 9735 24157
rect 9766 24148 9772 24200
rect 9824 24148 9830 24200
rect 9858 24148 9864 24200
rect 9916 24188 9922 24200
rect 10045 24191 10103 24197
rect 10045 24188 10057 24191
rect 9916 24160 10057 24188
rect 9916 24148 9922 24160
rect 10045 24157 10057 24160
rect 10091 24157 10103 24191
rect 10045 24151 10103 24157
rect 10321 24191 10379 24197
rect 10321 24157 10333 24191
rect 10367 24157 10379 24191
rect 10321 24151 10379 24157
rect 8987 24092 9352 24120
rect 9508 24120 9536 24148
rect 10336 24120 10364 24151
rect 10410 24148 10416 24200
rect 10468 24148 10474 24200
rect 9508 24092 10364 24120
rect 8987 24089 8999 24092
rect 8941 24083 8999 24089
rect 11790 24080 11796 24132
rect 11848 24080 11854 24132
rect 12066 24129 12072 24132
rect 12009 24123 12072 24129
rect 12009 24089 12021 24123
rect 12055 24089 12072 24123
rect 12009 24083 12072 24089
rect 12066 24080 12072 24083
rect 12124 24080 12130 24132
rect 12176 24120 12204 24228
rect 13725 24225 13737 24259
rect 13771 24256 13783 24259
rect 13771 24228 14228 24256
rect 13771 24225 13783 24228
rect 13725 24219 13783 24225
rect 12342 24148 12348 24200
rect 12400 24188 12406 24200
rect 12621 24191 12679 24197
rect 12621 24188 12633 24191
rect 12400 24160 12633 24188
rect 12400 24148 12406 24160
rect 12621 24157 12633 24160
rect 12667 24157 12679 24191
rect 12621 24151 12679 24157
rect 12710 24148 12716 24200
rect 12768 24188 12774 24200
rect 12897 24191 12955 24197
rect 12897 24188 12909 24191
rect 12768 24160 12909 24188
rect 12768 24148 12774 24160
rect 12897 24157 12909 24160
rect 12943 24157 12955 24191
rect 12897 24151 12955 24157
rect 12986 24148 12992 24200
rect 13044 24148 13050 24200
rect 13354 24148 13360 24200
rect 13412 24148 13418 24200
rect 14090 24148 14096 24200
rect 14148 24148 14154 24200
rect 14108 24120 14136 24148
rect 12176 24092 14136 24120
rect 14200 24120 14228 24228
rect 14292 24197 14320 24296
rect 17310 24284 17316 24336
rect 17368 24324 17374 24336
rect 17954 24324 17960 24336
rect 17368 24296 17960 24324
rect 17368 24284 17374 24296
rect 17954 24284 17960 24296
rect 18012 24284 18018 24336
rect 18064 24296 19288 24324
rect 15289 24259 15347 24265
rect 15289 24225 15301 24259
rect 15335 24256 15347 24259
rect 18064 24256 18092 24296
rect 19260 24268 19288 24296
rect 15335 24228 18092 24256
rect 15335 24225 15347 24228
rect 15289 24219 15347 24225
rect 18138 24216 18144 24268
rect 18196 24256 18202 24268
rect 19058 24256 19064 24268
rect 18196 24228 19064 24256
rect 18196 24216 18202 24228
rect 19058 24216 19064 24228
rect 19116 24216 19122 24268
rect 19242 24216 19248 24268
rect 19300 24216 19306 24268
rect 21836 24265 21864 24352
rect 23216 24324 23244 24364
rect 23290 24352 23296 24404
rect 23348 24392 23354 24404
rect 23845 24395 23903 24401
rect 23845 24392 23857 24395
rect 23348 24364 23857 24392
rect 23348 24352 23354 24364
rect 23845 24361 23857 24364
rect 23891 24361 23903 24395
rect 23845 24355 23903 24361
rect 24029 24395 24087 24401
rect 24029 24361 24041 24395
rect 24075 24392 24087 24395
rect 24946 24392 24952 24404
rect 24075 24364 24952 24392
rect 24075 24361 24087 24364
rect 24029 24355 24087 24361
rect 24946 24352 24952 24364
rect 25004 24352 25010 24404
rect 26326 24352 26332 24404
rect 26384 24352 26390 24404
rect 26421 24395 26479 24401
rect 26421 24361 26433 24395
rect 26467 24361 26479 24395
rect 27249 24395 27307 24401
rect 27249 24392 27261 24395
rect 26421 24355 26479 24361
rect 26988 24364 27261 24392
rect 24397 24327 24455 24333
rect 24397 24324 24409 24327
rect 23216 24296 24409 24324
rect 24397 24293 24409 24296
rect 24443 24293 24455 24327
rect 24397 24287 24455 24293
rect 25148 24296 25728 24324
rect 21821 24259 21879 24265
rect 21821 24225 21833 24259
rect 21867 24225 21879 24259
rect 21821 24219 21879 24225
rect 21910 24216 21916 24268
rect 21968 24216 21974 24268
rect 22554 24216 22560 24268
rect 22612 24256 22618 24268
rect 22612 24228 24256 24256
rect 22612 24216 22618 24228
rect 14277 24191 14335 24197
rect 14277 24157 14289 24191
rect 14323 24157 14335 24191
rect 14277 24151 14335 24157
rect 17218 24148 17224 24200
rect 17276 24198 17282 24200
rect 17276 24197 17356 24198
rect 17586 24197 17592 24200
rect 17276 24191 17371 24197
rect 17276 24170 17325 24191
rect 17276 24148 17282 24170
rect 17313 24157 17325 24170
rect 17359 24157 17371 24191
rect 17313 24151 17371 24157
rect 17543 24191 17592 24197
rect 17543 24157 17555 24191
rect 17589 24157 17592 24191
rect 17543 24151 17592 24157
rect 17586 24148 17592 24151
rect 17644 24148 17650 24200
rect 17678 24148 17684 24200
rect 17736 24148 17742 24200
rect 17770 24148 17776 24200
rect 17828 24148 17834 24200
rect 18233 24191 18291 24197
rect 18233 24157 18245 24191
rect 18279 24188 18291 24191
rect 18598 24188 18604 24200
rect 18279 24160 18604 24188
rect 18279 24157 18291 24160
rect 18233 24151 18291 24157
rect 18598 24148 18604 24160
rect 18656 24148 18662 24200
rect 20622 24148 20628 24200
rect 20680 24148 20686 24200
rect 21542 24148 21548 24200
rect 21600 24148 21606 24200
rect 14550 24120 14556 24132
rect 14200 24092 14556 24120
rect 14550 24080 14556 24092
rect 14608 24080 14614 24132
rect 15562 24080 15568 24132
rect 15620 24080 15626 24132
rect 16942 24120 16948 24132
rect 16790 24092 16948 24120
rect 16942 24080 16948 24092
rect 17000 24080 17006 24132
rect 17405 24123 17463 24129
rect 17405 24089 17417 24123
rect 17451 24120 17463 24123
rect 17451 24092 17908 24120
rect 17451 24089 17463 24092
rect 17405 24083 17463 24089
rect 17880 24064 17908 24092
rect 18966 24080 18972 24132
rect 19024 24120 19030 24132
rect 19521 24123 19579 24129
rect 19521 24120 19533 24123
rect 19024 24092 19533 24120
rect 19024 24080 19030 24092
rect 19521 24089 19533 24092
rect 19567 24089 19579 24123
rect 19521 24083 19579 24089
rect 20824 24092 22094 24120
rect 1578 24012 1584 24064
rect 1636 24012 1642 24064
rect 5169 24055 5227 24061
rect 5169 24021 5181 24055
rect 5215 24052 5227 24055
rect 5258 24052 5264 24064
rect 5215 24024 5264 24052
rect 5215 24021 5227 24024
rect 5169 24015 5227 24021
rect 5258 24012 5264 24024
rect 5316 24012 5322 24064
rect 14461 24055 14519 24061
rect 14461 24021 14473 24055
rect 14507 24052 14519 24055
rect 16206 24052 16212 24064
rect 14507 24024 16212 24052
rect 14507 24021 14519 24024
rect 14461 24015 14519 24021
rect 16206 24012 16212 24024
rect 16264 24052 16270 24064
rect 16482 24052 16488 24064
rect 16264 24024 16488 24052
rect 16264 24012 16270 24024
rect 16482 24012 16488 24024
rect 16540 24012 16546 24064
rect 16574 24012 16580 24064
rect 16632 24052 16638 24064
rect 17037 24055 17095 24061
rect 17037 24052 17049 24055
rect 16632 24024 17049 24052
rect 16632 24012 16638 24024
rect 17037 24021 17049 24024
rect 17083 24021 17095 24055
rect 17037 24015 17095 24021
rect 17126 24012 17132 24064
rect 17184 24012 17190 24064
rect 17862 24012 17868 24064
rect 17920 24012 17926 24064
rect 18046 24012 18052 24064
rect 18104 24052 18110 24064
rect 20824 24052 20852 24092
rect 18104 24024 20852 24052
rect 21361 24055 21419 24061
rect 18104 24012 18110 24024
rect 21361 24021 21373 24055
rect 21407 24052 21419 24055
rect 21818 24052 21824 24064
rect 21407 24024 21824 24052
rect 21407 24021 21419 24024
rect 21361 24015 21419 24021
rect 21818 24012 21824 24024
rect 21876 24012 21882 24064
rect 22066 24052 22094 24092
rect 22186 24080 22192 24132
rect 22244 24080 22250 24132
rect 23474 24120 23480 24132
rect 23414 24092 23480 24120
rect 23474 24080 23480 24092
rect 23532 24080 23538 24132
rect 24013 24123 24071 24129
rect 24013 24089 24025 24123
rect 24059 24120 24071 24123
rect 24118 24120 24124 24132
rect 24059 24092 24124 24120
rect 24059 24089 24071 24092
rect 24013 24083 24071 24089
rect 24118 24080 24124 24092
rect 24176 24080 24182 24132
rect 24228 24129 24256 24228
rect 24946 24216 24952 24268
rect 25004 24216 25010 24268
rect 25148 24265 25176 24296
rect 25133 24259 25191 24265
rect 25133 24225 25145 24259
rect 25179 24225 25191 24259
rect 25133 24219 25191 24225
rect 25498 24216 25504 24268
rect 25556 24256 25562 24268
rect 25593 24259 25651 24265
rect 25593 24256 25605 24259
rect 25556 24228 25605 24256
rect 25556 24216 25562 24228
rect 25593 24225 25605 24228
rect 25639 24225 25651 24259
rect 25700 24256 25728 24296
rect 25866 24284 25872 24336
rect 25924 24324 25930 24336
rect 26436 24324 26464 24355
rect 25924 24296 26464 24324
rect 25924 24284 25930 24296
rect 26988 24265 27016 24364
rect 27249 24361 27261 24364
rect 27295 24361 27307 24395
rect 27249 24355 27307 24361
rect 27433 24327 27491 24333
rect 27433 24293 27445 24327
rect 27479 24293 27491 24327
rect 27433 24287 27491 24293
rect 26973 24259 27031 24265
rect 26973 24256 26985 24259
rect 25700 24228 26985 24256
rect 25593 24219 25651 24225
rect 24302 24148 24308 24200
rect 24360 24188 24366 24200
rect 24670 24188 24676 24200
rect 24360 24160 24676 24188
rect 24360 24148 24366 24160
rect 24670 24148 24676 24160
rect 24728 24148 24734 24200
rect 25225 24191 25283 24197
rect 25225 24188 25237 24191
rect 24964 24160 25237 24188
rect 24213 24123 24271 24129
rect 24213 24089 24225 24123
rect 24259 24120 24271 24123
rect 24397 24123 24455 24129
rect 24397 24120 24409 24123
rect 24259 24092 24409 24120
rect 24259 24089 24271 24092
rect 24213 24083 24271 24089
rect 24397 24089 24409 24092
rect 24443 24089 24455 24123
rect 24762 24120 24768 24132
rect 24397 24083 24455 24089
rect 24504 24092 24768 24120
rect 23492 24052 23520 24080
rect 22066 24024 23520 24052
rect 23658 24012 23664 24064
rect 23716 24052 23722 24064
rect 24504 24052 24532 24092
rect 24762 24080 24768 24092
rect 24820 24120 24826 24132
rect 24964 24120 24992 24160
rect 25225 24157 25237 24160
rect 25271 24157 25283 24191
rect 25225 24151 25283 24157
rect 25682 24148 25688 24200
rect 25740 24148 25746 24200
rect 25866 24197 25872 24200
rect 25833 24191 25872 24197
rect 25833 24157 25845 24191
rect 25833 24151 25872 24157
rect 25866 24148 25872 24151
rect 25924 24148 25930 24200
rect 26068 24132 26096 24228
rect 26973 24225 26985 24228
rect 27019 24225 27031 24259
rect 26973 24219 27031 24225
rect 26142 24148 26148 24200
rect 26200 24197 26206 24200
rect 26200 24191 26249 24197
rect 26200 24157 26203 24191
rect 26237 24188 26249 24191
rect 26237 24160 26464 24188
rect 26237 24157 26249 24160
rect 26200 24151 26249 24157
rect 26200 24148 26206 24151
rect 24820 24092 24992 24120
rect 24820 24080 24826 24092
rect 25314 24080 25320 24132
rect 25372 24120 25378 24132
rect 25372 24092 25452 24120
rect 25372 24080 25378 24092
rect 23716 24024 24532 24052
rect 23716 24012 23722 24024
rect 24578 24012 24584 24064
rect 24636 24012 24642 24064
rect 25424 24061 25452 24092
rect 25498 24080 25504 24132
rect 25556 24080 25562 24132
rect 25590 24080 25596 24132
rect 25648 24120 25654 24132
rect 25961 24123 26019 24129
rect 25961 24120 25973 24123
rect 25648 24092 25973 24120
rect 25648 24080 25654 24092
rect 25961 24089 25973 24092
rect 26007 24089 26019 24123
rect 25961 24083 26019 24089
rect 26050 24080 26056 24132
rect 26108 24080 26114 24132
rect 26436 24120 26464 24160
rect 26510 24148 26516 24200
rect 26568 24188 26574 24200
rect 26605 24191 26663 24197
rect 26605 24188 26617 24191
rect 26568 24160 26617 24188
rect 26568 24148 26574 24160
rect 26605 24157 26617 24160
rect 26651 24157 26663 24191
rect 27448 24188 27476 24287
rect 27525 24191 27583 24197
rect 27525 24188 27537 24191
rect 27448 24160 27537 24188
rect 26605 24151 26663 24157
rect 27525 24157 27537 24160
rect 27571 24157 27583 24191
rect 27525 24151 27583 24157
rect 26436 24092 26832 24120
rect 26804 24061 26832 24092
rect 26878 24080 26884 24132
rect 26936 24120 26942 24132
rect 27065 24123 27123 24129
rect 27065 24120 27077 24123
rect 26936 24092 27077 24120
rect 26936 24080 26942 24092
rect 27065 24089 27077 24092
rect 27111 24089 27123 24123
rect 27065 24083 27123 24089
rect 27154 24080 27160 24132
rect 27212 24120 27218 24132
rect 27265 24123 27323 24129
rect 27265 24120 27277 24123
rect 27212 24092 27277 24120
rect 27212 24080 27218 24092
rect 27265 24089 27277 24092
rect 27311 24089 27323 24123
rect 27265 24083 27323 24089
rect 25409 24055 25467 24061
rect 25409 24021 25421 24055
rect 25455 24021 25467 24055
rect 25409 24015 25467 24021
rect 26789 24055 26847 24061
rect 26789 24021 26801 24055
rect 26835 24021 26847 24055
rect 26789 24015 26847 24021
rect 27706 24012 27712 24064
rect 27764 24012 27770 24064
rect 1104 23962 28152 23984
rect 1104 23910 4874 23962
rect 4926 23910 4938 23962
rect 4990 23910 5002 23962
rect 5054 23910 5066 23962
rect 5118 23910 5130 23962
rect 5182 23910 28152 23962
rect 1104 23888 28152 23910
rect 1578 23808 1584 23860
rect 1636 23848 1642 23860
rect 1636 23820 3372 23848
rect 1636 23808 1642 23820
rect 3050 23780 3056 23792
rect 2424 23752 3056 23780
rect 1486 23672 1492 23724
rect 1544 23672 1550 23724
rect 2424 23721 2452 23752
rect 3050 23740 3056 23752
rect 3108 23780 3114 23792
rect 3145 23783 3203 23789
rect 3145 23780 3157 23783
rect 3108 23752 3157 23780
rect 3108 23740 3114 23752
rect 3145 23749 3157 23752
rect 3191 23749 3203 23783
rect 3145 23743 3203 23749
rect 2409 23715 2467 23721
rect 2409 23681 2421 23715
rect 2455 23681 2467 23715
rect 2409 23675 2467 23681
rect 2498 23672 2504 23724
rect 2556 23672 2562 23724
rect 3344 23712 3372 23820
rect 3418 23808 3424 23860
rect 3476 23848 3482 23860
rect 8941 23851 8999 23857
rect 3476 23820 5488 23848
rect 3476 23808 3482 23820
rect 5350 23780 5356 23792
rect 5276 23752 5356 23780
rect 3513 23715 3571 23721
rect 3513 23712 3525 23715
rect 3344 23684 3525 23712
rect 3513 23681 3525 23684
rect 3559 23681 3571 23715
rect 3513 23675 3571 23681
rect 4341 23715 4399 23721
rect 4341 23681 4353 23715
rect 4387 23712 4399 23715
rect 4614 23712 4620 23724
rect 4387 23684 4620 23712
rect 4387 23681 4399 23684
rect 4341 23675 4399 23681
rect 3050 23604 3056 23656
rect 3108 23604 3114 23656
rect 2774 23536 2780 23588
rect 2832 23576 2838 23588
rect 3418 23576 3424 23588
rect 2832 23548 3424 23576
rect 2832 23536 2838 23548
rect 3418 23536 3424 23548
rect 3476 23536 3482 23588
rect 3528 23576 3556 23675
rect 4614 23672 4620 23684
rect 4672 23672 4678 23724
rect 4706 23672 4712 23724
rect 4764 23712 4770 23724
rect 5276 23721 5304 23752
rect 5350 23740 5356 23752
rect 5408 23740 5414 23792
rect 5261 23715 5319 23721
rect 4764 23684 5212 23712
rect 4764 23672 4770 23684
rect 4430 23604 4436 23656
rect 4488 23604 4494 23656
rect 4798 23604 4804 23656
rect 4856 23644 4862 23656
rect 5184 23653 5212 23684
rect 5261 23681 5273 23715
rect 5307 23681 5319 23715
rect 5261 23675 5319 23681
rect 4893 23647 4951 23653
rect 4893 23644 4905 23647
rect 4856 23616 4905 23644
rect 4856 23604 4862 23616
rect 4893 23613 4905 23616
rect 4939 23613 4951 23647
rect 4893 23607 4951 23613
rect 5169 23647 5227 23653
rect 5169 23613 5181 23647
rect 5215 23613 5227 23647
rect 5460 23644 5488 23820
rect 8941 23817 8953 23851
rect 8987 23848 8999 23851
rect 9861 23851 9919 23857
rect 8987 23820 9536 23848
rect 8987 23817 8999 23820
rect 8941 23811 8999 23817
rect 8570 23740 8576 23792
rect 8628 23780 8634 23792
rect 9508 23789 9536 23820
rect 9861 23817 9873 23851
rect 9907 23848 9919 23851
rect 10410 23848 10416 23860
rect 9907 23820 10416 23848
rect 9907 23817 9919 23820
rect 9861 23811 9919 23817
rect 10410 23808 10416 23820
rect 10468 23808 10474 23860
rect 12434 23848 12440 23860
rect 12084 23820 12440 23848
rect 9493 23783 9551 23789
rect 8628 23752 9076 23780
rect 8628 23740 8634 23752
rect 8846 23672 8852 23724
rect 8904 23672 8910 23724
rect 9048 23721 9076 23752
rect 9493 23749 9505 23783
rect 9539 23780 9551 23783
rect 9766 23780 9772 23792
rect 9539 23752 9772 23780
rect 9539 23749 9551 23752
rect 9493 23743 9551 23749
rect 9766 23740 9772 23752
rect 9824 23740 9830 23792
rect 9033 23715 9091 23721
rect 9033 23681 9045 23715
rect 9079 23681 9091 23715
rect 9033 23675 9091 23681
rect 9398 23672 9404 23724
rect 9456 23712 9462 23724
rect 12084 23721 12112 23820
rect 12434 23808 12440 23820
rect 12492 23808 12498 23860
rect 16390 23808 16396 23860
rect 16448 23848 16454 23860
rect 16853 23851 16911 23857
rect 16853 23848 16865 23851
rect 16448 23820 16865 23848
rect 16448 23808 16454 23820
rect 16853 23817 16865 23820
rect 16899 23817 16911 23851
rect 16853 23811 16911 23817
rect 17310 23808 17316 23860
rect 17368 23848 17374 23860
rect 17497 23851 17555 23857
rect 17497 23848 17509 23851
rect 17368 23820 17509 23848
rect 17368 23808 17374 23820
rect 17497 23817 17509 23820
rect 17543 23817 17555 23851
rect 17497 23811 17555 23817
rect 17589 23851 17647 23857
rect 17589 23817 17601 23851
rect 17635 23848 17647 23851
rect 17862 23848 17868 23860
rect 17635 23820 17868 23848
rect 17635 23817 17647 23820
rect 17589 23811 17647 23817
rect 17862 23808 17868 23820
rect 17920 23848 17926 23860
rect 17973 23851 18031 23857
rect 17973 23848 17985 23851
rect 17920 23820 17985 23848
rect 17920 23808 17926 23820
rect 17973 23817 17985 23820
rect 18019 23817 18031 23851
rect 17973 23811 18031 23817
rect 18966 23808 18972 23860
rect 19024 23808 19030 23860
rect 21542 23808 21548 23860
rect 21600 23848 21606 23860
rect 23753 23851 23811 23857
rect 23753 23848 23765 23851
rect 21600 23820 23765 23848
rect 21600 23808 21606 23820
rect 23753 23817 23765 23820
rect 23799 23817 23811 23851
rect 23753 23811 23811 23817
rect 24946 23808 24952 23860
rect 25004 23848 25010 23860
rect 25409 23851 25467 23857
rect 25409 23848 25421 23851
rect 25004 23820 25421 23848
rect 25004 23808 25010 23820
rect 25409 23817 25421 23820
rect 25455 23817 25467 23851
rect 25409 23811 25467 23817
rect 25866 23808 25872 23860
rect 25924 23848 25930 23860
rect 26878 23848 26884 23860
rect 25924 23820 26884 23848
rect 25924 23808 25930 23820
rect 26878 23808 26884 23820
rect 26936 23808 26942 23860
rect 13354 23780 13360 23792
rect 12820 23752 13360 23780
rect 9677 23715 9735 23721
rect 9677 23712 9689 23715
rect 9456 23684 9689 23712
rect 9456 23672 9462 23684
rect 9677 23681 9689 23684
rect 9723 23681 9735 23715
rect 9677 23675 9735 23681
rect 12069 23715 12127 23721
rect 12069 23681 12081 23715
rect 12115 23681 12127 23715
rect 12069 23675 12127 23681
rect 12250 23672 12256 23724
rect 12308 23672 12314 23724
rect 12434 23672 12440 23724
rect 12492 23672 12498 23724
rect 12621 23715 12679 23721
rect 12621 23681 12633 23715
rect 12667 23712 12679 23715
rect 12820 23712 12848 23752
rect 13354 23740 13360 23752
rect 13412 23740 13418 23792
rect 16761 23783 16819 23789
rect 16761 23780 16773 23783
rect 15948 23752 16773 23780
rect 15948 23724 15976 23752
rect 16761 23749 16773 23752
rect 16807 23749 16819 23783
rect 17402 23780 17408 23792
rect 16761 23743 16819 23749
rect 17144 23752 17408 23780
rect 12667 23684 12848 23712
rect 13173 23715 13231 23721
rect 12667 23681 12679 23684
rect 12621 23675 12679 23681
rect 13173 23681 13185 23715
rect 13219 23712 13231 23715
rect 14550 23712 14556 23724
rect 13219 23684 14556 23712
rect 13219 23681 13231 23684
rect 13173 23675 13231 23681
rect 14550 23672 14556 23684
rect 14608 23672 14614 23724
rect 15746 23672 15752 23724
rect 15804 23672 15810 23724
rect 15930 23672 15936 23724
rect 15988 23672 15994 23724
rect 16485 23715 16543 23721
rect 16485 23681 16497 23715
rect 16531 23712 16543 23715
rect 16574 23712 16580 23724
rect 16531 23684 16580 23712
rect 16531 23681 16543 23684
rect 16485 23675 16543 23681
rect 16574 23672 16580 23684
rect 16632 23672 16638 23724
rect 17144 23721 17172 23752
rect 17402 23740 17408 23752
rect 17460 23740 17466 23792
rect 17773 23783 17831 23789
rect 17773 23780 17785 23783
rect 17512 23752 17785 23780
rect 17512 23724 17540 23752
rect 17773 23749 17785 23752
rect 17819 23749 17831 23783
rect 17773 23743 17831 23749
rect 22002 23740 22008 23792
rect 22060 23780 22066 23792
rect 22097 23783 22155 23789
rect 22097 23780 22109 23783
rect 22060 23752 22109 23780
rect 22060 23740 22066 23752
rect 22097 23749 22109 23752
rect 22143 23749 22155 23783
rect 23474 23780 23480 23792
rect 23322 23752 23480 23780
rect 22097 23743 22155 23749
rect 23474 23740 23480 23752
rect 23532 23780 23538 23792
rect 25130 23780 25136 23792
rect 23532 23752 25136 23780
rect 23532 23740 23538 23752
rect 25130 23740 25136 23752
rect 25188 23740 25194 23792
rect 25314 23740 25320 23792
rect 25372 23780 25378 23792
rect 25501 23783 25559 23789
rect 25501 23780 25513 23783
rect 25372 23752 25513 23780
rect 25372 23740 25378 23752
rect 25501 23749 25513 23752
rect 25547 23749 25559 23783
rect 25501 23743 25559 23749
rect 16669 23715 16727 23721
rect 16669 23681 16681 23715
rect 16715 23681 16727 23715
rect 16669 23675 16727 23681
rect 17129 23715 17187 23721
rect 17129 23681 17141 23715
rect 17175 23681 17187 23715
rect 17129 23675 17187 23681
rect 17313 23715 17371 23721
rect 17313 23681 17325 23715
rect 17359 23712 17371 23715
rect 17494 23712 17500 23724
rect 17359 23684 17500 23712
rect 17359 23681 17371 23684
rect 17313 23675 17371 23681
rect 5460 23616 11284 23644
rect 5169 23607 5227 23613
rect 10318 23576 10324 23588
rect 3528 23548 10324 23576
rect 10318 23536 10324 23548
rect 10376 23536 10382 23588
rect 11256 23576 11284 23616
rect 12158 23604 12164 23656
rect 12216 23644 12222 23656
rect 12345 23647 12403 23653
rect 12345 23644 12357 23647
rect 12216 23616 12357 23644
rect 12216 23604 12222 23616
rect 12345 23613 12357 23616
rect 12391 23613 12403 23647
rect 12345 23607 12403 23613
rect 12897 23647 12955 23653
rect 12897 23613 12909 23647
rect 12943 23613 12955 23647
rect 15764 23644 15792 23672
rect 16684 23644 16712 23675
rect 17494 23672 17500 23684
rect 17552 23672 17558 23724
rect 17681 23715 17739 23721
rect 17681 23681 17693 23715
rect 17727 23712 17739 23715
rect 17862 23712 17868 23724
rect 17727 23684 17868 23712
rect 17727 23681 17739 23684
rect 17681 23675 17739 23681
rect 17862 23672 17868 23684
rect 17920 23672 17926 23724
rect 18598 23672 18604 23724
rect 18656 23672 18662 23724
rect 18874 23672 18880 23724
rect 18932 23672 18938 23724
rect 19426 23672 19432 23724
rect 19484 23672 19490 23724
rect 19610 23672 19616 23724
rect 19668 23672 19674 23724
rect 19705 23715 19763 23721
rect 19705 23681 19717 23715
rect 19751 23712 19763 23715
rect 20438 23712 20444 23724
rect 19751 23684 20444 23712
rect 19751 23681 19763 23684
rect 19705 23675 19763 23681
rect 20438 23672 20444 23684
rect 20496 23672 20502 23724
rect 21726 23672 21732 23724
rect 21784 23712 21790 23724
rect 21821 23715 21879 23721
rect 21821 23712 21833 23715
rect 21784 23684 21833 23712
rect 21784 23672 21790 23684
rect 21821 23681 21833 23684
rect 21867 23681 21879 23715
rect 21821 23675 21879 23681
rect 15764 23616 16712 23644
rect 12897 23607 12955 23613
rect 12912 23576 12940 23607
rect 17218 23604 17224 23656
rect 17276 23644 17282 23656
rect 19245 23647 19303 23653
rect 19245 23644 19257 23647
rect 17276 23616 19257 23644
rect 17276 23604 17282 23616
rect 19245 23613 19257 23616
rect 19291 23613 19303 23647
rect 19245 23607 19303 23613
rect 11256 23548 12940 23576
rect 17129 23579 17187 23585
rect 17129 23545 17141 23579
rect 17175 23576 17187 23579
rect 17678 23576 17684 23588
rect 17175 23548 17684 23576
rect 17175 23545 17187 23548
rect 17129 23539 17187 23545
rect 17678 23536 17684 23548
rect 17736 23536 17742 23588
rect 18506 23576 18512 23588
rect 17880 23548 18512 23576
rect 1765 23511 1823 23517
rect 1765 23477 1777 23511
rect 1811 23508 1823 23511
rect 2038 23508 2044 23520
rect 1811 23480 2044 23508
rect 1811 23477 1823 23480
rect 1765 23471 1823 23477
rect 2038 23468 2044 23480
rect 2096 23468 2102 23520
rect 5626 23468 5632 23520
rect 5684 23468 5690 23520
rect 12158 23468 12164 23520
rect 12216 23468 12222 23520
rect 12805 23511 12863 23517
rect 12805 23477 12817 23511
rect 12851 23508 12863 23511
rect 12986 23508 12992 23520
rect 12851 23480 12992 23508
rect 12851 23477 12863 23480
rect 12805 23471 12863 23477
rect 12986 23468 12992 23480
rect 13044 23468 13050 23520
rect 13357 23511 13415 23517
rect 13357 23477 13369 23511
rect 13403 23508 13415 23511
rect 15378 23508 15384 23520
rect 13403 23480 15384 23508
rect 13403 23477 13415 23480
rect 13357 23471 13415 23477
rect 15378 23468 15384 23480
rect 15436 23468 15442 23520
rect 15841 23511 15899 23517
rect 15841 23477 15853 23511
rect 15887 23508 15899 23511
rect 15930 23508 15936 23520
rect 15887 23480 15936 23508
rect 15887 23477 15899 23480
rect 15841 23471 15899 23477
rect 15930 23468 15936 23480
rect 15988 23508 15994 23520
rect 16298 23508 16304 23520
rect 15988 23480 16304 23508
rect 15988 23468 15994 23480
rect 16298 23468 16304 23480
rect 16356 23468 16362 23520
rect 16390 23468 16396 23520
rect 16448 23468 16454 23520
rect 16482 23468 16488 23520
rect 16540 23508 16546 23520
rect 17037 23511 17095 23517
rect 17037 23508 17049 23511
rect 16540 23480 17049 23508
rect 16540 23468 16546 23480
rect 17037 23477 17049 23480
rect 17083 23477 17095 23511
rect 17037 23471 17095 23477
rect 17405 23511 17463 23517
rect 17405 23477 17417 23511
rect 17451 23508 17463 23511
rect 17494 23508 17500 23520
rect 17451 23480 17500 23508
rect 17451 23477 17463 23480
rect 17405 23471 17463 23477
rect 17494 23468 17500 23480
rect 17552 23468 17558 23520
rect 17586 23468 17592 23520
rect 17644 23508 17650 23520
rect 17880 23508 17908 23548
rect 18506 23536 18512 23548
rect 18564 23576 18570 23588
rect 18693 23579 18751 23585
rect 18693 23576 18705 23579
rect 18564 23548 18705 23576
rect 18564 23536 18570 23548
rect 18693 23545 18705 23548
rect 18739 23545 18751 23579
rect 18693 23539 18751 23545
rect 17644 23480 17908 23508
rect 17644 23468 17650 23480
rect 17954 23468 17960 23520
rect 18012 23468 18018 23520
rect 18046 23468 18052 23520
rect 18104 23508 18110 23520
rect 18141 23511 18199 23517
rect 18141 23508 18153 23511
rect 18104 23480 18153 23508
rect 18104 23468 18110 23480
rect 18141 23477 18153 23480
rect 18187 23477 18199 23511
rect 21836 23508 21864 23675
rect 23382 23672 23388 23724
rect 23440 23712 23446 23724
rect 23661 23715 23719 23721
rect 23661 23712 23673 23715
rect 23440 23684 23673 23712
rect 23440 23672 23446 23684
rect 23661 23681 23673 23684
rect 23707 23681 23719 23715
rect 23661 23675 23719 23681
rect 23845 23715 23903 23721
rect 23845 23681 23857 23715
rect 23891 23712 23903 23715
rect 24026 23712 24032 23724
rect 23891 23684 24032 23712
rect 23891 23681 23903 23684
rect 23845 23675 23903 23681
rect 23106 23604 23112 23656
rect 23164 23644 23170 23656
rect 23860 23644 23888 23675
rect 24026 23672 24032 23684
rect 24084 23672 24090 23724
rect 24949 23715 25007 23721
rect 24949 23681 24961 23715
rect 24995 23712 25007 23715
rect 25590 23712 25596 23724
rect 24995 23684 25596 23712
rect 24995 23681 25007 23684
rect 24949 23675 25007 23681
rect 25590 23672 25596 23684
rect 25648 23672 25654 23724
rect 25685 23715 25743 23721
rect 25685 23681 25697 23715
rect 25731 23681 25743 23715
rect 25685 23675 25743 23681
rect 23164 23616 23888 23644
rect 23164 23604 23170 23616
rect 25038 23604 25044 23656
rect 25096 23644 25102 23656
rect 25498 23644 25504 23656
rect 25096 23616 25504 23644
rect 25096 23604 25102 23616
rect 25498 23604 25504 23616
rect 25556 23604 25562 23656
rect 23566 23536 23572 23588
rect 23624 23576 23630 23588
rect 25700 23576 25728 23675
rect 27522 23672 27528 23724
rect 27580 23672 27586 23724
rect 23624 23548 25728 23576
rect 23624 23536 23630 23548
rect 23474 23508 23480 23520
rect 21836 23480 23480 23508
rect 18141 23471 18199 23477
rect 23474 23468 23480 23480
rect 23532 23468 23538 23520
rect 24210 23468 24216 23520
rect 24268 23508 24274 23520
rect 24765 23511 24823 23517
rect 24765 23508 24777 23511
rect 24268 23480 24777 23508
rect 24268 23468 24274 23480
rect 24765 23477 24777 23480
rect 24811 23477 24823 23511
rect 24765 23471 24823 23477
rect 27706 23468 27712 23520
rect 27764 23468 27770 23520
rect 1104 23418 28152 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 28152 23418
rect 1104 23344 28152 23366
rect 4341 23307 4399 23313
rect 4341 23273 4353 23307
rect 4387 23304 4399 23307
rect 4614 23304 4620 23316
rect 4387 23276 4620 23304
rect 4387 23273 4399 23276
rect 4341 23267 4399 23273
rect 4614 23264 4620 23276
rect 4672 23264 4678 23316
rect 10413 23307 10471 23313
rect 10413 23273 10425 23307
rect 10459 23304 10471 23307
rect 11790 23304 11796 23316
rect 10459 23276 11796 23304
rect 10459 23273 10471 23276
rect 10413 23267 10471 23273
rect 11790 23264 11796 23276
rect 11848 23264 11854 23316
rect 12986 23264 12992 23316
rect 13044 23264 13050 23316
rect 19061 23307 19119 23313
rect 19061 23273 19073 23307
rect 19107 23304 19119 23307
rect 19610 23304 19616 23316
rect 19107 23276 19616 23304
rect 19107 23273 19119 23276
rect 19061 23267 19119 23273
rect 19610 23264 19616 23276
rect 19668 23264 19674 23316
rect 22186 23264 22192 23316
rect 22244 23304 22250 23316
rect 22465 23307 22523 23313
rect 22465 23304 22477 23307
rect 22244 23276 22477 23304
rect 22244 23264 22250 23276
rect 22465 23273 22477 23276
rect 22511 23273 22523 23307
rect 22465 23267 22523 23273
rect 22833 23307 22891 23313
rect 22833 23273 22845 23307
rect 22879 23304 22891 23307
rect 23382 23304 23388 23316
rect 22879 23276 23388 23304
rect 22879 23273 22891 23276
rect 22833 23267 22891 23273
rect 23382 23264 23388 23276
rect 23440 23264 23446 23316
rect 26789 23307 26847 23313
rect 26789 23273 26801 23307
rect 26835 23304 26847 23307
rect 27522 23304 27528 23316
rect 26835 23276 27528 23304
rect 26835 23273 26847 23276
rect 26789 23267 26847 23273
rect 27522 23264 27528 23276
rect 27580 23264 27586 23316
rect 4893 23239 4951 23245
rect 4893 23205 4905 23239
rect 4939 23236 4951 23239
rect 8205 23239 8263 23245
rect 4939 23208 5580 23236
rect 4939 23205 4951 23208
rect 4893 23199 4951 23205
rect 5552 23180 5580 23208
rect 8205 23205 8217 23239
rect 8251 23236 8263 23239
rect 8846 23236 8852 23248
rect 8251 23208 8852 23236
rect 8251 23205 8263 23208
rect 8205 23199 8263 23205
rect 8846 23196 8852 23208
rect 8904 23196 8910 23248
rect 9306 23196 9312 23248
rect 9364 23236 9370 23248
rect 10965 23239 11023 23245
rect 9364 23208 10824 23236
rect 9364 23196 9370 23208
rect 5169 23171 5227 23177
rect 4264 23140 5120 23168
rect 4264 23109 4292 23140
rect 4249 23103 4307 23109
rect 4249 23069 4261 23103
rect 4295 23069 4307 23103
rect 4249 23063 4307 23069
rect 4433 23103 4491 23109
rect 4433 23069 4445 23103
rect 4479 23100 4491 23103
rect 4614 23100 4620 23112
rect 4479 23072 4620 23100
rect 4479 23069 4491 23072
rect 4433 23063 4491 23069
rect 4614 23060 4620 23072
rect 4672 23060 4678 23112
rect 4706 23060 4712 23112
rect 4764 23100 4770 23112
rect 5092 23109 5120 23140
rect 5169 23137 5181 23171
rect 5215 23168 5227 23171
rect 5258 23168 5264 23180
rect 5215 23140 5264 23168
rect 5215 23137 5227 23140
rect 5169 23131 5227 23137
rect 5258 23128 5264 23140
rect 5316 23128 5322 23180
rect 5534 23128 5540 23180
rect 5592 23128 5598 23180
rect 7282 23128 7288 23180
rect 7340 23168 7346 23180
rect 7377 23171 7435 23177
rect 7377 23168 7389 23171
rect 7340 23140 7389 23168
rect 7340 23128 7346 23140
rect 7377 23137 7389 23140
rect 7423 23137 7435 23171
rect 7377 23131 7435 23137
rect 9217 23171 9275 23177
rect 9217 23137 9229 23171
rect 9263 23168 9275 23171
rect 10318 23168 10324 23180
rect 9263 23140 10324 23168
rect 9263 23137 9275 23140
rect 9217 23131 9275 23137
rect 10318 23128 10324 23140
rect 10376 23168 10382 23180
rect 10376 23140 10640 23168
rect 10376 23128 10382 23140
rect 6276 23112 6328 23118
rect 4893 23103 4951 23109
rect 4893 23100 4905 23103
rect 4764 23072 4905 23100
rect 4764 23060 4770 23072
rect 4893 23069 4905 23072
rect 4939 23069 4951 23103
rect 4893 23063 4951 23069
rect 5077 23103 5135 23109
rect 5077 23069 5089 23103
rect 5123 23100 5135 23103
rect 5442 23100 5448 23112
rect 5123 23072 5448 23100
rect 5123 23069 5135 23072
rect 5077 23063 5135 23069
rect 5442 23060 5448 23072
rect 5500 23060 5506 23112
rect 5626 23060 5632 23112
rect 5684 23060 5690 23112
rect 5813 23103 5871 23109
rect 5813 23069 5825 23103
rect 5859 23100 5871 23103
rect 6178 23100 6184 23112
rect 5859 23072 6184 23100
rect 5859 23069 5871 23072
rect 5813 23063 5871 23069
rect 6178 23060 6184 23072
rect 6236 23060 6242 23112
rect 7466 23060 7472 23112
rect 7524 23060 7530 23112
rect 7926 23060 7932 23112
rect 7984 23060 7990 23112
rect 8846 23060 8852 23112
rect 8904 23100 8910 23112
rect 9125 23103 9183 23109
rect 9125 23100 9137 23103
rect 8904 23072 9137 23100
rect 8904 23060 8910 23072
rect 9125 23069 9137 23072
rect 9171 23069 9183 23103
rect 9125 23063 9183 23069
rect 9306 23060 9312 23112
rect 9364 23100 9370 23112
rect 9401 23103 9459 23109
rect 9401 23100 9413 23103
rect 9364 23072 9413 23100
rect 9364 23060 9370 23072
rect 9401 23069 9413 23072
rect 9447 23069 9459 23103
rect 9401 23063 9459 23069
rect 9490 23060 9496 23112
rect 9548 23100 9554 23112
rect 9769 23103 9827 23109
rect 9548 23072 9720 23100
rect 9548 23060 9554 23072
rect 6276 23054 6328 23060
rect 7193 23035 7251 23041
rect 7193 23001 7205 23035
rect 7239 23032 7251 23035
rect 7282 23032 7288 23044
rect 7239 23004 7288 23032
rect 7239 23001 7251 23004
rect 7193 22995 7251 23001
rect 7282 22992 7288 23004
rect 7340 22992 7346 23044
rect 8205 23035 8263 23041
rect 8205 23032 8217 23035
rect 7852 23004 8217 23032
rect 7852 22976 7880 23004
rect 8205 23001 8217 23004
rect 8251 23001 8263 23035
rect 8205 22995 8263 23001
rect 9585 23035 9643 23041
rect 9585 23001 9597 23035
rect 9631 23001 9643 23035
rect 9692 23032 9720 23072
rect 9769 23069 9781 23103
rect 9815 23100 9827 23103
rect 9861 23103 9919 23109
rect 9861 23100 9873 23103
rect 9815 23072 9873 23100
rect 9815 23069 9827 23072
rect 9769 23063 9827 23069
rect 9861 23069 9873 23072
rect 9907 23069 9919 23103
rect 9861 23063 9919 23069
rect 9950 23060 9956 23112
rect 10008 23060 10014 23112
rect 10137 23103 10195 23109
rect 10137 23069 10149 23103
rect 10183 23069 10195 23103
rect 10137 23063 10195 23069
rect 10152 23032 10180 23063
rect 10226 23060 10232 23112
rect 10284 23060 10290 23112
rect 10502 23060 10508 23112
rect 10560 23060 10566 23112
rect 10612 23109 10640 23140
rect 10796 23109 10824 23208
rect 10965 23205 10977 23239
rect 11011 23236 11023 23239
rect 19334 23236 19340 23248
rect 11011 23208 19340 23236
rect 11011 23205 11023 23208
rect 10965 23199 11023 23205
rect 12805 23171 12863 23177
rect 12805 23137 12817 23171
rect 12851 23168 12863 23171
rect 14274 23168 14280 23180
rect 12851 23140 14280 23168
rect 12851 23137 12863 23140
rect 12805 23131 12863 23137
rect 14274 23128 14280 23140
rect 14332 23128 14338 23180
rect 10597 23103 10655 23109
rect 10597 23069 10609 23103
rect 10643 23069 10655 23103
rect 10597 23063 10655 23069
rect 10781 23103 10839 23109
rect 10781 23069 10793 23103
rect 10827 23069 10839 23103
rect 10781 23063 10839 23069
rect 12250 23060 12256 23112
rect 12308 23100 12314 23112
rect 12345 23103 12403 23109
rect 12345 23100 12357 23103
rect 12308 23072 12357 23100
rect 12308 23060 12314 23072
rect 12345 23069 12357 23072
rect 12391 23069 12403 23103
rect 12345 23063 12403 23069
rect 12437 23103 12495 23109
rect 12437 23069 12449 23103
rect 12483 23100 12495 23103
rect 12526 23100 12532 23112
rect 12483 23072 12532 23100
rect 12483 23069 12495 23072
rect 12437 23063 12495 23069
rect 9692 23004 10180 23032
rect 12360 23032 12388 23063
rect 12526 23060 12532 23072
rect 12584 23060 12590 23112
rect 12618 23060 12624 23112
rect 12676 23060 12682 23112
rect 12894 23060 12900 23112
rect 12952 23060 12958 23112
rect 13262 23060 13268 23112
rect 13320 23060 13326 23112
rect 13538 23060 13544 23112
rect 13596 23100 13602 23112
rect 18708 23109 18736 23208
rect 19334 23196 19340 23208
rect 19392 23196 19398 23248
rect 19426 23196 19432 23248
rect 19484 23236 19490 23248
rect 19981 23239 20039 23245
rect 19981 23236 19993 23239
rect 19484 23208 19993 23236
rect 19484 23196 19490 23208
rect 19981 23205 19993 23208
rect 20027 23236 20039 23239
rect 20349 23239 20407 23245
rect 20349 23236 20361 23239
rect 20027 23208 20361 23236
rect 20027 23205 20039 23208
rect 19981 23199 20039 23205
rect 20349 23205 20361 23208
rect 20395 23205 20407 23239
rect 23658 23236 23664 23248
rect 20349 23199 20407 23205
rect 22940 23208 23664 23236
rect 22940 23177 22968 23208
rect 23658 23196 23664 23208
rect 23716 23196 23722 23248
rect 26234 23196 26240 23248
rect 26292 23236 26298 23248
rect 26697 23239 26755 23245
rect 26697 23236 26709 23239
rect 26292 23208 26709 23236
rect 26292 23196 26298 23208
rect 26697 23205 26709 23208
rect 26743 23205 26755 23239
rect 26697 23199 26755 23205
rect 22925 23171 22983 23177
rect 19076 23140 20392 23168
rect 19076 23109 19104 23140
rect 20364 23112 20392 23140
rect 22925 23137 22937 23171
rect 22971 23137 22983 23171
rect 22925 23131 22983 23137
rect 23474 23128 23480 23180
rect 23532 23168 23538 23180
rect 24394 23168 24400 23180
rect 23532 23140 24400 23168
rect 23532 23128 23538 23140
rect 24394 23128 24400 23140
rect 24452 23128 24458 23180
rect 18509 23103 18567 23109
rect 18509 23100 18521 23103
rect 13596 23072 18521 23100
rect 13596 23060 13602 23072
rect 18509 23069 18521 23072
rect 18555 23069 18567 23103
rect 18509 23063 18567 23069
rect 18693 23103 18751 23109
rect 18693 23069 18705 23103
rect 18739 23100 18751 23103
rect 18969 23103 19027 23109
rect 18969 23100 18981 23103
rect 18739 23072 18981 23100
rect 18739 23069 18751 23072
rect 18693 23063 18751 23069
rect 18969 23069 18981 23072
rect 19015 23069 19027 23103
rect 18969 23063 19027 23069
rect 19061 23103 19119 23109
rect 19061 23069 19073 23103
rect 19107 23069 19119 23103
rect 20073 23103 20131 23109
rect 20073 23100 20085 23103
rect 19061 23063 19119 23069
rect 19260 23072 20085 23100
rect 12912 23032 12940 23060
rect 12360 23004 12940 23032
rect 18524 23032 18552 23063
rect 18785 23035 18843 23041
rect 18785 23032 18797 23035
rect 18524 23004 18797 23032
rect 9585 22995 9643 23001
rect 18785 23001 18797 23004
rect 18831 23001 18843 23035
rect 18785 22995 18843 23001
rect 4614 22924 4620 22976
rect 4672 22964 4678 22976
rect 4890 22964 4896 22976
rect 4672 22936 4896 22964
rect 4672 22924 4678 22936
rect 4890 22924 4896 22936
rect 4948 22924 4954 22976
rect 7834 22924 7840 22976
rect 7892 22924 7898 22976
rect 8018 22924 8024 22976
rect 8076 22924 8082 22976
rect 9600 22964 9628 22995
rect 9766 22964 9772 22976
rect 9600 22936 9772 22964
rect 9766 22924 9772 22936
rect 9824 22924 9830 22976
rect 13449 22967 13507 22973
rect 13449 22933 13461 22967
rect 13495 22964 13507 22967
rect 14090 22964 14096 22976
rect 13495 22936 14096 22964
rect 13495 22933 13507 22936
rect 13449 22927 13507 22933
rect 14090 22924 14096 22936
rect 14148 22924 14154 22976
rect 18690 22924 18696 22976
rect 18748 22924 18754 22976
rect 18800 22964 18828 22995
rect 19260 22964 19288 23072
rect 20073 23069 20085 23072
rect 20119 23069 20131 23103
rect 20073 23063 20131 23069
rect 20346 23060 20352 23112
rect 20404 23060 20410 23112
rect 20438 23060 20444 23112
rect 20496 23060 20502 23112
rect 20625 23103 20683 23109
rect 20625 23069 20637 23103
rect 20671 23100 20683 23103
rect 20806 23100 20812 23112
rect 20671 23072 20812 23100
rect 20671 23069 20683 23072
rect 20625 23063 20683 23069
rect 20806 23060 20812 23072
rect 20864 23060 20870 23112
rect 22649 23103 22707 23109
rect 22649 23069 22661 23103
rect 22695 23100 22707 23103
rect 22738 23100 22744 23112
rect 22695 23072 22744 23100
rect 22695 23069 22707 23072
rect 22649 23063 22707 23069
rect 22738 23060 22744 23072
rect 22796 23060 22802 23112
rect 23201 23103 23259 23109
rect 23201 23069 23213 23103
rect 23247 23100 23259 23103
rect 23842 23100 23848 23112
rect 23247 23072 23848 23100
rect 23247 23069 23259 23072
rect 23201 23063 23259 23069
rect 23842 23060 23848 23072
rect 23900 23060 23906 23112
rect 24026 23060 24032 23112
rect 24084 23060 24090 23112
rect 24210 23060 24216 23112
rect 24268 23060 24274 23112
rect 26142 23060 26148 23112
rect 26200 23100 26206 23112
rect 26605 23103 26663 23109
rect 26605 23100 26617 23103
rect 26200 23072 26617 23100
rect 26200 23060 26206 23072
rect 26605 23069 26617 23072
rect 26651 23069 26663 23103
rect 26605 23063 26663 23069
rect 19334 22992 19340 23044
rect 19392 23032 19398 23044
rect 19613 23035 19671 23041
rect 19392 23004 19564 23032
rect 19392 22992 19398 23004
rect 18800 22936 19288 22964
rect 19426 22924 19432 22976
rect 19484 22924 19490 22976
rect 19536 22964 19564 23004
rect 19613 23001 19625 23035
rect 19659 23032 19671 23035
rect 19659 23004 20300 23032
rect 19659 23001 19671 23004
rect 19613 22995 19671 23001
rect 20165 22967 20223 22973
rect 20165 22964 20177 22967
rect 19536 22936 20177 22964
rect 20165 22933 20177 22936
rect 20211 22933 20223 22967
rect 20272 22964 20300 23004
rect 22462 22992 22468 23044
rect 22520 23032 22526 23044
rect 23017 23035 23075 23041
rect 23017 23032 23029 23035
rect 22520 23004 23029 23032
rect 22520 22992 22526 23004
rect 23017 23001 23029 23004
rect 23063 23001 23075 23035
rect 23017 22995 23075 23001
rect 20533 22967 20591 22973
rect 20533 22964 20545 22967
rect 20272 22936 20545 22964
rect 20165 22927 20223 22933
rect 20533 22933 20545 22936
rect 20579 22933 20591 22967
rect 24044 22964 24072 23060
rect 24121 23035 24179 23041
rect 24121 23001 24133 23035
rect 24167 23032 24179 23035
rect 24673 23035 24731 23041
rect 24673 23032 24685 23035
rect 24167 23004 24685 23032
rect 24167 23001 24179 23004
rect 24121 22995 24179 23001
rect 24673 23001 24685 23004
rect 24719 23001 24731 23035
rect 24673 22995 24731 23001
rect 25130 22992 25136 23044
rect 25188 22992 25194 23044
rect 26878 22992 26884 23044
rect 26936 22992 26942 23044
rect 25498 22964 25504 22976
rect 24044 22936 25504 22964
rect 20533 22927 20591 22933
rect 25498 22924 25504 22936
rect 25556 22924 25562 22976
rect 25958 22924 25964 22976
rect 26016 22964 26022 22976
rect 26145 22967 26203 22973
rect 26145 22964 26157 22967
rect 26016 22936 26157 22964
rect 26016 22924 26022 22936
rect 26145 22933 26157 22936
rect 26191 22933 26203 22967
rect 26145 22927 26203 22933
rect 1104 22874 28152 22896
rect 1104 22822 4874 22874
rect 4926 22822 4938 22874
rect 4990 22822 5002 22874
rect 5054 22822 5066 22874
rect 5118 22822 5130 22874
rect 5182 22822 28152 22874
rect 1104 22800 28152 22822
rect 3142 22760 3148 22772
rect 2424 22732 3148 22760
rect 842 22652 848 22704
rect 900 22692 906 22704
rect 1489 22695 1547 22701
rect 1489 22692 1501 22695
rect 900 22664 1501 22692
rect 900 22652 906 22664
rect 1489 22661 1501 22664
rect 1535 22661 1547 22695
rect 1489 22655 1547 22661
rect 2222 22584 2228 22636
rect 2280 22584 2286 22636
rect 2424 22633 2452 22732
rect 3142 22720 3148 22732
rect 3200 22720 3206 22772
rect 7834 22720 7840 22772
rect 7892 22760 7898 22772
rect 7945 22763 8003 22769
rect 7945 22760 7957 22763
rect 7892 22732 7957 22760
rect 7892 22720 7898 22732
rect 7945 22729 7957 22732
rect 7991 22729 8003 22763
rect 7945 22723 8003 22729
rect 8113 22763 8171 22769
rect 8113 22729 8125 22763
rect 8159 22760 8171 22763
rect 10226 22760 10232 22772
rect 8159 22732 8708 22760
rect 8159 22729 8171 22732
rect 8113 22723 8171 22729
rect 8680 22701 8708 22732
rect 9692 22732 10232 22760
rect 6549 22695 6607 22701
rect 3068 22664 3924 22692
rect 3068 22636 3096 22664
rect 2409 22627 2467 22633
rect 2409 22593 2421 22627
rect 2455 22593 2467 22627
rect 2409 22587 2467 22593
rect 3050 22584 3056 22636
rect 3108 22584 3114 22636
rect 3896 22633 3924 22664
rect 6549 22661 6561 22695
rect 6595 22692 6607 22695
rect 7745 22695 7803 22701
rect 7745 22692 7757 22695
rect 6595 22664 7757 22692
rect 6595 22661 6607 22664
rect 6549 22655 6607 22661
rect 7745 22661 7757 22664
rect 7791 22692 7803 22695
rect 8665 22695 8723 22701
rect 7791 22664 8064 22692
rect 7791 22661 7803 22664
rect 7745 22655 7803 22661
rect 8036 22636 8064 22664
rect 8665 22661 8677 22695
rect 8711 22661 8723 22695
rect 8665 22655 8723 22661
rect 8846 22652 8852 22704
rect 8904 22652 8910 22704
rect 9398 22652 9404 22704
rect 9456 22692 9462 22704
rect 9585 22695 9643 22701
rect 9585 22692 9597 22695
rect 9456 22664 9597 22692
rect 9456 22652 9462 22664
rect 9585 22661 9597 22664
rect 9631 22661 9643 22695
rect 9585 22655 9643 22661
rect 3697 22627 3755 22633
rect 3697 22593 3709 22627
rect 3743 22593 3755 22627
rect 3697 22587 3755 22593
rect 3881 22627 3939 22633
rect 3881 22593 3893 22627
rect 3927 22593 3939 22627
rect 3881 22587 3939 22593
rect 2317 22559 2375 22565
rect 2317 22525 2329 22559
rect 2363 22556 2375 22559
rect 2777 22559 2835 22565
rect 2777 22556 2789 22559
rect 2363 22528 2789 22556
rect 2363 22525 2375 22528
rect 2317 22519 2375 22525
rect 2777 22525 2789 22528
rect 2823 22556 2835 22559
rect 2823 22528 3096 22556
rect 2823 22525 2835 22528
rect 2777 22519 2835 22525
rect 1673 22491 1731 22497
rect 1673 22457 1685 22491
rect 1719 22488 1731 22491
rect 3068 22488 3096 22528
rect 3602 22516 3608 22568
rect 3660 22516 3666 22568
rect 3712 22488 3740 22587
rect 5534 22584 5540 22636
rect 5592 22584 5598 22636
rect 6178 22584 6184 22636
rect 6236 22624 6242 22636
rect 6457 22627 6515 22633
rect 6457 22624 6469 22627
rect 6236 22596 6469 22624
rect 6236 22584 6242 22596
rect 6457 22593 6469 22596
rect 6503 22593 6515 22627
rect 6457 22587 6515 22593
rect 6641 22627 6699 22633
rect 6641 22593 6653 22627
rect 6687 22593 6699 22627
rect 6641 22587 6699 22593
rect 5626 22516 5632 22568
rect 5684 22516 5690 22568
rect 6270 22516 6276 22568
rect 6328 22556 6334 22568
rect 6656 22556 6684 22587
rect 8018 22584 8024 22636
rect 8076 22584 8082 22636
rect 9214 22584 9220 22636
rect 9272 22624 9278 22636
rect 9493 22627 9551 22633
rect 9493 22624 9505 22627
rect 9272 22596 9505 22624
rect 9272 22584 9278 22596
rect 9493 22593 9505 22596
rect 9539 22624 9551 22627
rect 9692 22624 9720 22732
rect 10226 22720 10232 22732
rect 10284 22720 10290 22772
rect 10321 22763 10379 22769
rect 10321 22729 10333 22763
rect 10367 22760 10379 22763
rect 13538 22760 13544 22772
rect 10367 22732 13544 22760
rect 10367 22729 10379 22732
rect 10321 22723 10379 22729
rect 13538 22720 13544 22732
rect 13596 22720 13602 22772
rect 13633 22763 13691 22769
rect 13633 22729 13645 22763
rect 13679 22760 13691 22763
rect 14293 22763 14351 22769
rect 14293 22760 14305 22763
rect 13679 22732 14305 22760
rect 13679 22729 13691 22732
rect 13633 22723 13691 22729
rect 14293 22729 14305 22732
rect 14339 22729 14351 22763
rect 14293 22723 14351 22729
rect 17129 22763 17187 22769
rect 17129 22729 17141 22763
rect 17175 22760 17187 22763
rect 17310 22760 17316 22772
rect 17175 22732 17316 22760
rect 17175 22729 17187 22732
rect 17129 22723 17187 22729
rect 17310 22720 17316 22732
rect 17368 22720 17374 22772
rect 17862 22720 17868 22772
rect 17920 22760 17926 22772
rect 19426 22760 19432 22772
rect 17920 22732 19432 22760
rect 17920 22720 17926 22732
rect 19426 22720 19432 22732
rect 19484 22720 19490 22772
rect 20806 22720 20812 22772
rect 20864 22720 20870 22772
rect 26418 22720 26424 22772
rect 26476 22760 26482 22772
rect 27173 22763 27231 22769
rect 27173 22760 27185 22763
rect 26476 22732 27185 22760
rect 26476 22720 26482 22732
rect 27173 22729 27185 22732
rect 27219 22729 27231 22763
rect 27173 22723 27231 22729
rect 9858 22652 9864 22704
rect 9916 22692 9922 22704
rect 9953 22695 10011 22701
rect 9953 22692 9965 22695
rect 9916 22664 9965 22692
rect 9916 22652 9922 22664
rect 9953 22661 9965 22664
rect 9999 22692 10011 22695
rect 10502 22692 10508 22704
rect 9999 22664 10508 22692
rect 9999 22661 10011 22664
rect 9953 22655 10011 22661
rect 9539 22596 9720 22624
rect 9539 22593 9551 22596
rect 9493 22587 9551 22593
rect 9766 22584 9772 22636
rect 9824 22584 9830 22636
rect 10042 22584 10048 22636
rect 10100 22584 10106 22636
rect 10244 22633 10272 22664
rect 10502 22652 10508 22664
rect 10560 22652 10566 22704
rect 14090 22652 14096 22704
rect 14148 22652 14154 22704
rect 16574 22652 16580 22704
rect 16632 22692 16638 22704
rect 16761 22695 16819 22701
rect 16761 22692 16773 22695
rect 16632 22664 16773 22692
rect 16632 22652 16638 22664
rect 16761 22661 16773 22664
rect 16807 22661 16819 22695
rect 16761 22655 16819 22661
rect 16977 22695 17035 22701
rect 16977 22661 16989 22695
rect 17023 22692 17035 22695
rect 17023 22664 19472 22692
rect 17023 22661 17035 22664
rect 16977 22655 17035 22661
rect 10229 22627 10287 22633
rect 10229 22593 10241 22627
rect 10275 22593 10287 22627
rect 10229 22587 10287 22593
rect 10318 22584 10324 22636
rect 10376 22584 10382 22636
rect 12805 22627 12863 22633
rect 12805 22593 12817 22627
rect 12851 22593 12863 22627
rect 12805 22587 12863 22593
rect 13265 22627 13323 22633
rect 13265 22593 13277 22627
rect 13311 22624 13323 22627
rect 13354 22624 13360 22636
rect 13311 22596 13360 22624
rect 13311 22593 13323 22596
rect 13265 22587 13323 22593
rect 6328 22528 6684 22556
rect 9033 22559 9091 22565
rect 6328 22516 6334 22528
rect 9033 22525 9045 22559
rect 9079 22556 9091 22559
rect 9784 22556 9812 22584
rect 9079 22528 9812 22556
rect 9079 22525 9091 22528
rect 9033 22519 9091 22525
rect 12710 22488 12716 22500
rect 1719 22460 3004 22488
rect 3068 22460 3740 22488
rect 3804 22460 12716 22488
rect 1719 22457 1731 22460
rect 1673 22451 1731 22457
rect 2130 22380 2136 22432
rect 2188 22420 2194 22432
rect 2406 22420 2412 22432
rect 2188 22392 2412 22420
rect 2188 22380 2194 22392
rect 2406 22380 2412 22392
rect 2464 22380 2470 22432
rect 2976 22420 3004 22460
rect 3234 22420 3240 22432
rect 2976 22392 3240 22420
rect 3234 22380 3240 22392
rect 3292 22420 3298 22432
rect 3804 22420 3832 22460
rect 12710 22448 12716 22460
rect 12768 22448 12774 22500
rect 12820 22488 12848 22587
rect 13354 22584 13360 22596
rect 13412 22584 13418 22636
rect 16776 22624 16804 22655
rect 17512 22633 17540 22664
rect 17221 22627 17279 22633
rect 17221 22624 17233 22627
rect 16776 22596 17233 22624
rect 17221 22593 17233 22596
rect 17267 22593 17279 22627
rect 17221 22587 17279 22593
rect 17405 22627 17463 22633
rect 17405 22593 17417 22627
rect 17451 22593 17463 22627
rect 17405 22587 17463 22593
rect 17497 22627 17555 22633
rect 17497 22593 17509 22627
rect 17543 22593 17555 22627
rect 18598 22624 18604 22636
rect 17497 22587 17555 22593
rect 17604 22596 18604 22624
rect 13078 22516 13084 22568
rect 13136 22556 13142 22568
rect 13173 22559 13231 22565
rect 13173 22556 13185 22559
rect 13136 22528 13185 22556
rect 13136 22516 13142 22528
rect 13173 22525 13185 22528
rect 13219 22556 13231 22559
rect 13722 22556 13728 22568
rect 13219 22528 13728 22556
rect 13219 22525 13231 22528
rect 13173 22519 13231 22525
rect 13722 22516 13728 22528
rect 13780 22516 13786 22568
rect 17420 22556 17448 22587
rect 17604 22556 17632 22596
rect 18598 22584 18604 22596
rect 18656 22624 18662 22636
rect 19337 22627 19395 22633
rect 19337 22624 19349 22627
rect 18656 22596 19349 22624
rect 18656 22584 18662 22596
rect 19337 22593 19349 22596
rect 19383 22593 19395 22627
rect 19337 22587 19395 22593
rect 19444 22565 19472 22664
rect 20438 22652 20444 22704
rect 20496 22692 20502 22704
rect 21361 22695 21419 22701
rect 21361 22692 21373 22695
rect 20496 22664 21373 22692
rect 20496 22652 20502 22664
rect 21361 22661 21373 22664
rect 21407 22661 21419 22695
rect 21361 22655 21419 22661
rect 26878 22652 26884 22704
rect 26936 22692 26942 22704
rect 26973 22695 27031 22701
rect 26973 22692 26985 22695
rect 26936 22664 26985 22692
rect 26936 22652 26942 22664
rect 26973 22661 26985 22664
rect 27019 22661 27031 22695
rect 26973 22655 27031 22661
rect 20990 22584 20996 22636
rect 21048 22624 21054 22636
rect 21269 22627 21327 22633
rect 21269 22624 21281 22627
rect 21048 22596 21281 22624
rect 21048 22584 21054 22596
rect 21269 22593 21281 22596
rect 21315 22593 21327 22627
rect 21269 22587 21327 22593
rect 21453 22627 21511 22633
rect 21453 22593 21465 22627
rect 21499 22624 21511 22627
rect 22278 22624 22284 22636
rect 21499 22596 22284 22624
rect 21499 22593 21511 22596
rect 21453 22587 21511 22593
rect 17420 22528 17632 22556
rect 19429 22559 19487 22565
rect 13262 22488 13268 22500
rect 12820 22460 13268 22488
rect 13262 22448 13268 22460
rect 13320 22448 13326 22500
rect 17420 22488 17448 22528
rect 19429 22525 19441 22559
rect 19475 22556 19487 22559
rect 20530 22556 20536 22568
rect 19475 22528 20536 22556
rect 19475 22525 19487 22528
rect 19429 22519 19487 22525
rect 20530 22516 20536 22528
rect 20588 22516 20594 22568
rect 21177 22559 21235 22565
rect 21177 22525 21189 22559
rect 21223 22556 21235 22559
rect 21468 22556 21496 22587
rect 22278 22584 22284 22596
rect 22336 22584 22342 22636
rect 25682 22584 25688 22636
rect 25740 22584 25746 22636
rect 25869 22627 25927 22633
rect 25869 22593 25881 22627
rect 25915 22624 25927 22627
rect 25958 22624 25964 22636
rect 25915 22596 25964 22624
rect 25915 22593 25927 22596
rect 25869 22587 25927 22593
rect 25958 22584 25964 22596
rect 26016 22584 26022 22636
rect 26053 22627 26111 22633
rect 26053 22593 26065 22627
rect 26099 22624 26111 22627
rect 26142 22624 26148 22636
rect 26099 22596 26148 22624
rect 26099 22593 26111 22596
rect 26053 22587 26111 22593
rect 26142 22584 26148 22596
rect 26200 22624 26206 22636
rect 26513 22627 26571 22633
rect 26513 22624 26525 22627
rect 26200 22596 26525 22624
rect 26200 22584 26206 22596
rect 26513 22593 26525 22596
rect 26559 22593 26571 22627
rect 27525 22627 27583 22633
rect 27525 22624 27537 22627
rect 26513 22587 26571 22593
rect 27356 22596 27537 22624
rect 21223 22528 21496 22556
rect 21223 22525 21235 22528
rect 21177 22519 21235 22525
rect 27356 22497 27384 22596
rect 27525 22593 27537 22596
rect 27571 22593 27583 22627
rect 27525 22587 27583 22593
rect 16960 22460 17448 22488
rect 27341 22491 27399 22497
rect 3292 22392 3832 22420
rect 3292 22380 3298 22392
rect 3878 22380 3884 22432
rect 3936 22380 3942 22432
rect 5905 22423 5963 22429
rect 5905 22389 5917 22423
rect 5951 22420 5963 22423
rect 6362 22420 6368 22432
rect 5951 22392 6368 22420
rect 5951 22389 5963 22392
rect 5905 22383 5963 22389
rect 6362 22380 6368 22392
rect 6420 22380 6426 22432
rect 7374 22380 7380 22432
rect 7432 22420 7438 22432
rect 7926 22420 7932 22432
rect 7432 22392 7932 22420
rect 7432 22380 7438 22392
rect 7926 22380 7932 22392
rect 7984 22380 7990 22432
rect 9306 22380 9312 22432
rect 9364 22420 9370 22432
rect 10042 22420 10048 22432
rect 9364 22392 10048 22420
rect 9364 22380 9370 22392
rect 10042 22380 10048 22392
rect 10100 22380 10106 22432
rect 12618 22380 12624 22432
rect 12676 22420 12682 22432
rect 12802 22420 12808 22432
rect 12676 22392 12808 22420
rect 12676 22380 12682 22392
rect 12802 22380 12808 22392
rect 12860 22420 12866 22432
rect 12897 22423 12955 22429
rect 12897 22420 12909 22423
rect 12860 22392 12909 22420
rect 12860 22380 12866 22392
rect 12897 22389 12909 22392
rect 12943 22389 12955 22423
rect 12897 22383 12955 22389
rect 14274 22380 14280 22432
rect 14332 22380 14338 22432
rect 14461 22423 14519 22429
rect 14461 22389 14473 22423
rect 14507 22420 14519 22423
rect 16114 22420 16120 22432
rect 14507 22392 16120 22420
rect 14507 22389 14519 22392
rect 14461 22383 14519 22389
rect 16114 22380 16120 22392
rect 16172 22380 16178 22432
rect 16960 22429 16988 22460
rect 27341 22457 27353 22491
rect 27387 22457 27399 22491
rect 27341 22451 27399 22457
rect 27706 22448 27712 22500
rect 27764 22448 27770 22500
rect 16945 22423 17003 22429
rect 16945 22389 16957 22423
rect 16991 22389 17003 22423
rect 16945 22383 17003 22389
rect 17218 22380 17224 22432
rect 17276 22380 17282 22432
rect 19610 22380 19616 22432
rect 19668 22380 19674 22432
rect 25406 22380 25412 22432
rect 25464 22420 25470 22432
rect 25501 22423 25559 22429
rect 25501 22420 25513 22423
rect 25464 22392 25513 22420
rect 25464 22380 25470 22392
rect 25501 22389 25513 22392
rect 25547 22389 25559 22423
rect 25501 22383 25559 22389
rect 25958 22380 25964 22432
rect 26016 22380 26022 22432
rect 26234 22380 26240 22432
rect 26292 22420 26298 22432
rect 27157 22423 27215 22429
rect 27157 22420 27169 22423
rect 26292 22392 27169 22420
rect 26292 22380 26298 22392
rect 27157 22389 27169 22392
rect 27203 22389 27215 22423
rect 27157 22383 27215 22389
rect 1104 22330 28152 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 28152 22330
rect 1104 22256 28152 22278
rect 3053 22219 3111 22225
rect 3053 22185 3065 22219
rect 3099 22216 3111 22219
rect 3142 22216 3148 22228
rect 3099 22188 3148 22216
rect 3099 22185 3111 22188
rect 3053 22179 3111 22185
rect 2222 22040 2228 22092
rect 2280 22040 2286 22092
rect 842 21972 848 22024
rect 900 22012 906 22024
rect 1397 22015 1455 22021
rect 1397 22012 1409 22015
rect 900 21984 1409 22012
rect 900 21972 906 21984
rect 1397 21981 1409 21984
rect 1443 21981 1455 22015
rect 1397 21975 1455 21981
rect 2133 22015 2191 22021
rect 2133 21981 2145 22015
rect 2179 22012 2191 22015
rect 3068 22012 3096 22179
rect 3142 22176 3148 22188
rect 3200 22176 3206 22228
rect 4525 22219 4583 22225
rect 4525 22185 4537 22219
rect 4571 22216 4583 22219
rect 4706 22216 4712 22228
rect 4571 22188 4712 22216
rect 4571 22185 4583 22188
rect 4525 22179 4583 22185
rect 4154 22108 4160 22160
rect 4212 22108 4218 22160
rect 3878 22040 3884 22092
rect 3936 22040 3942 22092
rect 3973 22083 4031 22089
rect 3973 22049 3985 22083
rect 4019 22080 4031 22083
rect 4172 22080 4200 22108
rect 4540 22080 4568 22179
rect 4706 22176 4712 22188
rect 4764 22176 4770 22228
rect 7374 22176 7380 22228
rect 7432 22176 7438 22228
rect 20990 22216 20996 22228
rect 12406 22188 20996 22216
rect 12406 22148 12434 22188
rect 20990 22176 20996 22188
rect 21048 22216 21054 22228
rect 21542 22216 21548 22228
rect 21048 22188 21548 22216
rect 21048 22176 21054 22188
rect 21542 22176 21548 22188
rect 21600 22176 21606 22228
rect 25777 22219 25835 22225
rect 25777 22185 25789 22219
rect 25823 22216 25835 22219
rect 26234 22216 26240 22228
rect 25823 22188 26240 22216
rect 25823 22185 25835 22188
rect 25777 22179 25835 22185
rect 26234 22176 26240 22188
rect 26292 22176 26298 22228
rect 16206 22148 16212 22160
rect 10612 22120 12434 22148
rect 15304 22120 16212 22148
rect 10612 22089 10640 22120
rect 4019 22052 4568 22080
rect 9309 22083 9367 22089
rect 4019 22049 4031 22052
rect 3973 22043 4031 22049
rect 9309 22049 9321 22083
rect 9355 22080 9367 22083
rect 9677 22083 9735 22089
rect 9677 22080 9689 22083
rect 9355 22052 9689 22080
rect 9355 22049 9367 22052
rect 9309 22043 9367 22049
rect 9677 22049 9689 22052
rect 9723 22049 9735 22083
rect 9677 22043 9735 22049
rect 10597 22083 10655 22089
rect 10597 22049 10609 22083
rect 10643 22049 10655 22083
rect 10597 22043 10655 22049
rect 14274 22040 14280 22092
rect 14332 22080 14338 22092
rect 14332 22052 14964 22080
rect 14332 22040 14338 22052
rect 2179 21984 3096 22012
rect 2179 21981 2191 21984
rect 2133 21975 2191 21981
rect 3234 21972 3240 22024
rect 3292 21972 3298 22024
rect 3694 21972 3700 22024
rect 3752 22012 3758 22024
rect 4065 22015 4123 22021
rect 4065 22012 4077 22015
rect 3752 21984 4077 22012
rect 3752 21972 3758 21984
rect 4065 21981 4077 21984
rect 4111 21981 4123 22015
rect 4065 21975 4123 21981
rect 4157 22015 4215 22021
rect 4157 21981 4169 22015
rect 4203 21981 4215 22015
rect 4433 22015 4491 22021
rect 4433 22012 4445 22015
rect 4157 21975 4215 21981
rect 4264 21984 4445 22012
rect 3602 21904 3608 21956
rect 3660 21944 3666 21956
rect 3970 21944 3976 21956
rect 3660 21916 3976 21944
rect 3660 21904 3666 21916
rect 3970 21904 3976 21916
rect 4028 21944 4034 21956
rect 4172 21944 4200 21975
rect 4028 21916 4200 21944
rect 4028 21904 4034 21916
rect 1581 21879 1639 21885
rect 1581 21845 1593 21879
rect 1627 21876 1639 21879
rect 2774 21876 2780 21888
rect 1627 21848 2780 21876
rect 1627 21845 1639 21848
rect 1581 21839 1639 21845
rect 2774 21836 2780 21848
rect 2832 21836 2838 21888
rect 2866 21836 2872 21888
rect 2924 21836 2930 21888
rect 3418 21836 3424 21888
rect 3476 21876 3482 21888
rect 4264 21876 4292 21984
rect 4433 21981 4445 21984
rect 4479 22012 4491 22015
rect 4706 22012 4712 22024
rect 4479 21984 4712 22012
rect 4479 21981 4491 21984
rect 4433 21975 4491 21981
rect 4706 21972 4712 21984
rect 4764 21972 4770 22024
rect 7282 21972 7288 22024
rect 7340 21972 7346 22024
rect 7374 21972 7380 22024
rect 7432 22012 7438 22024
rect 7469 22015 7527 22021
rect 7469 22012 7481 22015
rect 7432 21984 7481 22012
rect 7432 21972 7438 21984
rect 7469 21981 7481 21984
rect 7515 21981 7527 22015
rect 7469 21975 7527 21981
rect 9214 21972 9220 22024
rect 9272 21972 9278 22024
rect 9398 21972 9404 22024
rect 9456 21972 9462 22024
rect 9766 21972 9772 22024
rect 9824 21972 9830 22024
rect 12342 21972 12348 22024
rect 12400 22012 12406 22024
rect 13354 22012 13360 22024
rect 12400 21984 13360 22012
rect 12400 21972 12406 21984
rect 13354 21972 13360 21984
rect 13412 21972 13418 22024
rect 13722 21972 13728 22024
rect 13780 21972 13786 22024
rect 14458 21972 14464 22024
rect 14516 22012 14522 22024
rect 14936 22021 14964 22052
rect 15304 22021 15332 22120
rect 16206 22108 16212 22120
rect 16264 22148 16270 22160
rect 16301 22151 16359 22157
rect 16301 22148 16313 22151
rect 16264 22120 16313 22148
rect 16264 22108 16270 22120
rect 16301 22117 16313 22120
rect 16347 22117 16359 22151
rect 26142 22148 26148 22160
rect 16301 22111 16359 22117
rect 25240 22120 26148 22148
rect 16853 22083 16911 22089
rect 16853 22049 16865 22083
rect 16899 22080 16911 22083
rect 17034 22080 17040 22092
rect 16899 22052 17040 22080
rect 16899 22049 16911 22052
rect 16853 22043 16911 22049
rect 17034 22040 17040 22052
rect 17092 22040 17098 22092
rect 14645 22015 14703 22021
rect 14645 22012 14657 22015
rect 14516 21984 14657 22012
rect 14516 21972 14522 21984
rect 14645 21981 14657 21984
rect 14691 21981 14703 22015
rect 14645 21975 14703 21981
rect 14921 22015 14979 22021
rect 14921 21981 14933 22015
rect 14967 21981 14979 22015
rect 14921 21975 14979 21981
rect 15289 22015 15347 22021
rect 15289 21981 15301 22015
rect 15335 21981 15347 22015
rect 15289 21975 15347 21981
rect 15473 22015 15531 22021
rect 15473 21981 15485 22015
rect 15519 22012 15531 22015
rect 17129 22015 17187 22021
rect 15519 21984 16344 22012
rect 15519 21981 15531 21984
rect 15473 21975 15531 21981
rect 13740 21944 13768 21972
rect 16316 21956 16344 21984
rect 17129 21981 17141 22015
rect 17175 22012 17187 22015
rect 17218 22012 17224 22024
rect 17175 21984 17224 22012
rect 17175 21981 17187 21984
rect 17129 21975 17187 21981
rect 17218 21972 17224 21984
rect 17276 21972 17282 22024
rect 17310 21972 17316 22024
rect 17368 21972 17374 22024
rect 24670 21972 24676 22024
rect 24728 22012 24734 22024
rect 25240 22021 25268 22120
rect 26142 22108 26148 22120
rect 26200 22108 26206 22160
rect 25774 22040 25780 22092
rect 25832 22080 25838 22092
rect 26418 22080 26424 22092
rect 25832 22052 26424 22080
rect 25832 22040 25838 22052
rect 26418 22040 26424 22052
rect 26476 22040 26482 22092
rect 25225 22015 25283 22021
rect 25225 22012 25237 22015
rect 24728 21984 25237 22012
rect 24728 21972 24734 21984
rect 25225 21981 25237 21984
rect 25271 21981 25283 22015
rect 25225 21975 25283 21981
rect 25314 21972 25320 22024
rect 25372 21972 25378 22024
rect 25682 21972 25688 22024
rect 25740 22012 25746 22024
rect 25740 21984 26096 22012
rect 25740 21972 25746 21984
rect 26068 21956 26096 21984
rect 14274 21944 14280 21956
rect 13740 21916 14280 21944
rect 14274 21904 14280 21916
rect 14332 21904 14338 21956
rect 16298 21904 16304 21956
rect 16356 21904 16362 21956
rect 25498 21904 25504 21956
rect 25556 21904 25562 21956
rect 25961 21947 26019 21953
rect 25961 21913 25973 21947
rect 26007 21913 26019 21947
rect 25961 21907 26019 21913
rect 3476 21848 4292 21876
rect 4341 21879 4399 21885
rect 3476 21836 3482 21848
rect 4341 21845 4353 21879
rect 4387 21876 4399 21879
rect 4614 21876 4620 21888
rect 4387 21848 4620 21876
rect 4387 21845 4399 21848
rect 4341 21839 4399 21845
rect 4614 21836 4620 21848
rect 4672 21836 4678 21888
rect 13449 21879 13507 21885
rect 13449 21845 13461 21879
rect 13495 21876 13507 21879
rect 13538 21876 13544 21888
rect 13495 21848 13544 21876
rect 13495 21845 13507 21848
rect 13449 21839 13507 21845
rect 13538 21836 13544 21848
rect 13596 21876 13602 21888
rect 14366 21876 14372 21888
rect 13596 21848 14372 21876
rect 13596 21836 13602 21848
rect 14366 21836 14372 21848
rect 14424 21836 14430 21888
rect 15194 21836 15200 21888
rect 15252 21836 15258 21888
rect 16114 21836 16120 21888
rect 16172 21876 16178 21888
rect 16761 21879 16819 21885
rect 16761 21876 16773 21879
rect 16172 21848 16773 21876
rect 16172 21836 16178 21848
rect 16761 21845 16773 21848
rect 16807 21845 16819 21879
rect 16761 21839 16819 21845
rect 17037 21879 17095 21885
rect 17037 21845 17049 21879
rect 17083 21876 17095 21879
rect 17126 21876 17132 21888
rect 17083 21848 17132 21876
rect 17083 21845 17095 21848
rect 17037 21839 17095 21845
rect 17126 21836 17132 21848
rect 17184 21836 17190 21888
rect 17497 21879 17555 21885
rect 17497 21845 17509 21879
rect 17543 21876 17555 21879
rect 17678 21876 17684 21888
rect 17543 21848 17684 21876
rect 17543 21845 17555 21848
rect 17497 21839 17555 21845
rect 17678 21836 17684 21848
rect 17736 21836 17742 21888
rect 25038 21836 25044 21888
rect 25096 21876 25102 21888
rect 25225 21879 25283 21885
rect 25225 21876 25237 21879
rect 25096 21848 25237 21876
rect 25096 21836 25102 21848
rect 25225 21845 25237 21848
rect 25271 21845 25283 21879
rect 25225 21839 25283 21845
rect 25590 21836 25596 21888
rect 25648 21836 25654 21888
rect 25774 21885 25780 21888
rect 25761 21879 25780 21885
rect 25761 21845 25773 21879
rect 25761 21839 25780 21845
rect 25774 21836 25780 21839
rect 25832 21836 25838 21888
rect 25976 21876 26004 21907
rect 26050 21904 26056 21956
rect 26108 21944 26114 21956
rect 26145 21947 26203 21953
rect 26145 21944 26157 21947
rect 26108 21916 26157 21944
rect 26108 21904 26114 21916
rect 26145 21913 26157 21916
rect 26191 21913 26203 21947
rect 26145 21907 26203 21913
rect 26237 21879 26295 21885
rect 26237 21876 26249 21879
rect 25976 21848 26249 21876
rect 26237 21845 26249 21848
rect 26283 21876 26295 21879
rect 26970 21876 26976 21888
rect 26283 21848 26976 21876
rect 26283 21845 26295 21848
rect 26237 21839 26295 21845
rect 26970 21836 26976 21848
rect 27028 21836 27034 21888
rect 1104 21786 28152 21808
rect 1104 21734 4874 21786
rect 4926 21734 4938 21786
rect 4990 21734 5002 21786
rect 5054 21734 5066 21786
rect 5118 21734 5130 21786
rect 5182 21734 28152 21786
rect 1104 21712 28152 21734
rect 2222 21672 2228 21684
rect 1964 21644 2228 21672
rect 1964 21613 1992 21644
rect 2222 21632 2228 21644
rect 2280 21632 2286 21684
rect 4433 21675 4491 21681
rect 4433 21641 4445 21675
rect 4479 21672 4491 21675
rect 4706 21672 4712 21684
rect 4479 21644 4712 21672
rect 4479 21641 4491 21644
rect 4433 21635 4491 21641
rect 4706 21632 4712 21644
rect 4764 21632 4770 21684
rect 13078 21632 13084 21684
rect 13136 21672 13142 21684
rect 13136 21644 14412 21672
rect 13136 21632 13142 21644
rect 1949 21607 2007 21613
rect 1949 21573 1961 21607
rect 1995 21573 2007 21607
rect 1949 21567 2007 21573
rect 12713 21607 12771 21613
rect 12713 21573 12725 21607
rect 12759 21604 12771 21607
rect 13357 21607 13415 21613
rect 13357 21604 13369 21607
rect 12759 21576 13369 21604
rect 12759 21573 12771 21576
rect 12713 21567 12771 21573
rect 13357 21573 13369 21576
rect 13403 21573 13415 21607
rect 14384 21604 14412 21644
rect 14458 21632 14464 21684
rect 14516 21632 14522 21684
rect 19702 21672 19708 21684
rect 19306 21644 19708 21672
rect 19306 21604 19334 21644
rect 19702 21632 19708 21644
rect 19760 21672 19766 21684
rect 23290 21672 23296 21684
rect 19760 21644 23296 21672
rect 19760 21632 19766 21644
rect 23290 21632 23296 21644
rect 23348 21632 23354 21684
rect 24946 21632 24952 21684
rect 25004 21672 25010 21684
rect 25251 21675 25309 21681
rect 25251 21672 25263 21675
rect 25004 21644 25263 21672
rect 25004 21632 25010 21644
rect 25251 21641 25263 21644
rect 25297 21672 25309 21675
rect 25958 21672 25964 21684
rect 25297 21644 25964 21672
rect 25297 21641 25309 21644
rect 25251 21635 25309 21641
rect 25958 21632 25964 21644
rect 26016 21632 26022 21684
rect 26053 21675 26111 21681
rect 26053 21641 26065 21675
rect 26099 21672 26111 21675
rect 26142 21672 26148 21684
rect 26099 21644 26148 21672
rect 26099 21641 26111 21644
rect 26053 21635 26111 21641
rect 26142 21632 26148 21644
rect 26200 21632 26206 21684
rect 14384 21576 19334 21604
rect 13357 21567 13415 21573
rect 19978 21564 19984 21616
rect 20036 21604 20042 21616
rect 20346 21604 20352 21616
rect 20036 21576 20352 21604
rect 20036 21564 20042 21576
rect 20346 21564 20352 21576
rect 20404 21604 20410 21616
rect 20441 21607 20499 21613
rect 20441 21604 20453 21607
rect 20404 21576 20453 21604
rect 20404 21564 20410 21576
rect 20441 21573 20453 21576
rect 20487 21573 20499 21607
rect 20441 21567 20499 21573
rect 24673 21607 24731 21613
rect 24673 21573 24685 21607
rect 24719 21604 24731 21607
rect 25041 21607 25099 21613
rect 25041 21604 25053 21607
rect 24719 21576 25053 21604
rect 24719 21573 24731 21576
rect 24673 21567 24731 21573
rect 25041 21573 25053 21576
rect 25087 21604 25099 21607
rect 25406 21604 25412 21616
rect 25087 21576 25412 21604
rect 25087 21573 25099 21576
rect 25041 21567 25099 21573
rect 25406 21564 25412 21576
rect 25464 21564 25470 21616
rect 25593 21607 25651 21613
rect 25593 21573 25605 21607
rect 25639 21604 25651 21607
rect 26234 21604 26240 21616
rect 25639 21576 26240 21604
rect 25639 21573 25651 21576
rect 25593 21567 25651 21573
rect 26234 21564 26240 21576
rect 26292 21564 26298 21616
rect 2682 21536 2688 21548
rect 2622 21508 2688 21536
rect 2682 21496 2688 21508
rect 2740 21496 2746 21548
rect 3786 21496 3792 21548
rect 3844 21496 3850 21548
rect 3970 21496 3976 21548
rect 4028 21496 4034 21548
rect 4614 21496 4620 21548
rect 4672 21496 4678 21548
rect 4982 21496 4988 21548
rect 5040 21496 5046 21548
rect 7374 21496 7380 21548
rect 7432 21496 7438 21548
rect 12342 21496 12348 21548
rect 12400 21536 12406 21548
rect 12621 21539 12679 21545
rect 12621 21536 12633 21539
rect 12400 21508 12633 21536
rect 12400 21496 12406 21508
rect 12621 21505 12633 21508
rect 12667 21505 12679 21539
rect 12621 21499 12679 21505
rect 12805 21539 12863 21545
rect 12805 21505 12817 21539
rect 12851 21536 12863 21539
rect 12894 21536 12900 21548
rect 12851 21508 12900 21536
rect 12851 21505 12863 21508
rect 12805 21499 12863 21505
rect 2498 21428 2504 21480
rect 2556 21428 2562 21480
rect 5629 21471 5687 21477
rect 5629 21437 5641 21471
rect 5675 21468 5687 21471
rect 5718 21468 5724 21480
rect 5675 21440 5724 21468
rect 5675 21437 5687 21440
rect 5629 21431 5687 21437
rect 5718 21428 5724 21440
rect 5776 21428 5782 21480
rect 7282 21428 7288 21480
rect 7340 21428 7346 21480
rect 8110 21428 8116 21480
rect 8168 21428 8174 21480
rect 12636 21468 12664 21499
rect 12894 21496 12900 21508
rect 12952 21496 12958 21548
rect 13078 21496 13084 21548
rect 13136 21496 13142 21548
rect 13170 21496 13176 21548
rect 13228 21496 13234 21548
rect 13541 21539 13599 21545
rect 13541 21536 13553 21539
rect 13464 21508 13553 21536
rect 13464 21468 13492 21508
rect 13541 21505 13553 21508
rect 13587 21505 13599 21539
rect 13541 21499 13599 21505
rect 13630 21496 13636 21548
rect 13688 21534 13694 21548
rect 13909 21539 13967 21545
rect 13688 21506 13731 21534
rect 13688 21496 13694 21506
rect 13909 21505 13921 21539
rect 13955 21536 13967 21539
rect 14090 21536 14096 21548
rect 13955 21508 14096 21536
rect 13955 21505 13967 21508
rect 13909 21499 13967 21505
rect 14090 21496 14096 21508
rect 14148 21496 14154 21548
rect 14274 21496 14280 21548
rect 14332 21496 14338 21548
rect 14918 21496 14924 21548
rect 14976 21496 14982 21548
rect 15102 21496 15108 21548
rect 15160 21496 15166 21548
rect 16114 21496 16120 21548
rect 16172 21496 16178 21548
rect 16298 21496 16304 21548
rect 16356 21496 16362 21548
rect 17126 21496 17132 21548
rect 17184 21496 17190 21548
rect 17589 21539 17647 21545
rect 17589 21505 17601 21539
rect 17635 21505 17647 21539
rect 17589 21499 17647 21505
rect 12636 21440 13492 21468
rect 15289 21471 15347 21477
rect 15289 21437 15301 21471
rect 15335 21468 15347 21471
rect 16206 21468 16212 21480
rect 15335 21440 16212 21468
rect 15335 21437 15347 21440
rect 15289 21431 15347 21437
rect 16206 21428 16212 21440
rect 16264 21428 16270 21480
rect 16485 21471 16543 21477
rect 16485 21437 16497 21471
rect 16531 21468 16543 21471
rect 17402 21468 17408 21480
rect 16531 21440 17408 21468
rect 16531 21437 16543 21440
rect 16485 21431 16543 21437
rect 17402 21428 17408 21440
rect 17460 21468 17466 21480
rect 17604 21468 17632 21499
rect 18046 21496 18052 21548
rect 18104 21496 18110 21548
rect 18417 21539 18475 21545
rect 18417 21505 18429 21539
rect 18463 21505 18475 21539
rect 18417 21499 18475 21505
rect 18969 21539 19027 21545
rect 18969 21505 18981 21539
rect 19015 21505 19027 21539
rect 18969 21499 19027 21505
rect 17460 21440 17632 21468
rect 17460 21428 17466 21440
rect 17862 21428 17868 21480
rect 17920 21468 17926 21480
rect 18432 21468 18460 21499
rect 17920 21440 18460 21468
rect 18984 21468 19012 21499
rect 19058 21496 19064 21548
rect 19116 21536 19122 21548
rect 19613 21539 19671 21545
rect 19613 21536 19625 21539
rect 19116 21508 19625 21536
rect 19116 21496 19122 21508
rect 19613 21505 19625 21508
rect 19659 21505 19671 21539
rect 19613 21499 19671 21505
rect 20533 21539 20591 21545
rect 20533 21505 20545 21539
rect 20579 21536 20591 21539
rect 21082 21536 21088 21548
rect 20579 21508 21088 21536
rect 20579 21505 20591 21508
rect 20533 21499 20591 21505
rect 21082 21496 21088 21508
rect 21140 21496 21146 21548
rect 23106 21496 23112 21548
rect 23164 21496 23170 21548
rect 24857 21539 24915 21545
rect 24857 21505 24869 21539
rect 24903 21505 24915 21539
rect 24857 21499 24915 21505
rect 19426 21468 19432 21480
rect 18984 21440 19432 21468
rect 17920 21428 17926 21440
rect 12526 21360 12532 21412
rect 12584 21400 12590 21412
rect 13078 21400 13084 21412
rect 12584 21372 13084 21400
rect 12584 21360 12590 21372
rect 13078 21360 13084 21372
rect 13136 21360 13142 21412
rect 13170 21360 13176 21412
rect 13228 21400 13234 21412
rect 13722 21400 13728 21412
rect 13228 21372 13728 21400
rect 13228 21360 13234 21372
rect 13722 21360 13728 21372
rect 13780 21400 13786 21412
rect 13817 21403 13875 21409
rect 13817 21400 13829 21403
rect 13780 21372 13829 21400
rect 13780 21360 13786 21372
rect 13817 21369 13829 21372
rect 13863 21369 13875 21403
rect 14366 21400 14372 21412
rect 13817 21363 13875 21369
rect 14292 21372 14372 21400
rect 12897 21335 12955 21341
rect 12897 21301 12909 21335
rect 12943 21332 12955 21335
rect 12986 21332 12992 21344
rect 12943 21304 12992 21332
rect 12943 21301 12955 21304
rect 12897 21295 12955 21301
rect 12986 21292 12992 21304
rect 13044 21292 13050 21344
rect 13357 21335 13415 21341
rect 13357 21301 13369 21335
rect 13403 21332 13415 21335
rect 13630 21332 13636 21344
rect 13403 21304 13636 21332
rect 13403 21301 13415 21304
rect 13357 21295 13415 21301
rect 13630 21292 13636 21304
rect 13688 21292 13694 21344
rect 14292 21341 14320 21372
rect 14366 21360 14372 21372
rect 14424 21360 14430 21412
rect 17218 21360 17224 21412
rect 17276 21360 17282 21412
rect 17770 21360 17776 21412
rect 17828 21400 17834 21412
rect 18984 21400 19012 21440
rect 19426 21428 19432 21440
rect 19484 21428 19490 21480
rect 22186 21428 22192 21480
rect 22244 21468 22250 21480
rect 22922 21468 22928 21480
rect 22244 21440 22928 21468
rect 22244 21428 22250 21440
rect 22922 21428 22928 21440
rect 22980 21428 22986 21480
rect 24872 21468 24900 21499
rect 24946 21496 24952 21548
rect 25004 21496 25010 21548
rect 25501 21539 25559 21545
rect 25501 21505 25513 21539
rect 25547 21505 25559 21539
rect 25501 21499 25559 21505
rect 25130 21468 25136 21480
rect 24872 21440 25136 21468
rect 25130 21428 25136 21440
rect 25188 21428 25194 21480
rect 17828 21372 19012 21400
rect 17828 21360 17834 21372
rect 21174 21360 21180 21412
rect 21232 21400 21238 21412
rect 22738 21400 22744 21412
rect 21232 21372 22744 21400
rect 21232 21360 21238 21372
rect 22738 21360 22744 21372
rect 22796 21360 22802 21412
rect 24673 21403 24731 21409
rect 24673 21369 24685 21403
rect 24719 21400 24731 21403
rect 25314 21400 25320 21412
rect 24719 21372 25320 21400
rect 24719 21369 24731 21372
rect 24673 21363 24731 21369
rect 25314 21360 25320 21372
rect 25372 21360 25378 21412
rect 25409 21403 25467 21409
rect 25409 21369 25421 21403
rect 25455 21400 25467 21403
rect 25516 21400 25544 21499
rect 25682 21496 25688 21548
rect 25740 21536 25746 21548
rect 25777 21539 25835 21545
rect 25777 21536 25789 21539
rect 25740 21508 25789 21536
rect 25740 21496 25746 21508
rect 25777 21505 25789 21508
rect 25823 21505 25835 21539
rect 25777 21499 25835 21505
rect 27154 21496 27160 21548
rect 27212 21496 27218 21548
rect 25590 21428 25596 21480
rect 25648 21468 25654 21480
rect 26513 21471 26571 21477
rect 26513 21468 26525 21471
rect 25648 21440 26525 21468
rect 25648 21428 25654 21440
rect 26513 21437 26525 21440
rect 26559 21437 26571 21471
rect 26513 21431 26571 21437
rect 26142 21400 26148 21412
rect 25455 21372 26148 21400
rect 25455 21369 25467 21372
rect 25409 21363 25467 21369
rect 26142 21360 26148 21372
rect 26200 21360 26206 21412
rect 26970 21360 26976 21412
rect 27028 21360 27034 21412
rect 14277 21335 14335 21341
rect 14277 21301 14289 21335
rect 14323 21301 14335 21335
rect 14277 21295 14335 21301
rect 16022 21292 16028 21344
rect 16080 21332 16086 21344
rect 19518 21332 19524 21344
rect 16080 21304 19524 21332
rect 16080 21292 16086 21304
rect 19518 21292 19524 21304
rect 19576 21332 19582 21344
rect 19794 21332 19800 21344
rect 19576 21304 19800 21332
rect 19576 21292 19582 21304
rect 19794 21292 19800 21304
rect 19852 21292 19858 21344
rect 21358 21292 21364 21344
rect 21416 21332 21422 21344
rect 22833 21335 22891 21341
rect 22833 21332 22845 21335
rect 21416 21304 22845 21332
rect 21416 21292 21422 21304
rect 22833 21301 22845 21304
rect 22879 21332 22891 21335
rect 23014 21332 23020 21344
rect 22879 21304 23020 21332
rect 22879 21301 22891 21304
rect 22833 21295 22891 21301
rect 23014 21292 23020 21304
rect 23072 21292 23078 21344
rect 25130 21292 25136 21344
rect 25188 21332 25194 21344
rect 25225 21335 25283 21341
rect 25225 21332 25237 21335
rect 25188 21304 25237 21332
rect 25188 21292 25194 21304
rect 25225 21301 25237 21304
rect 25271 21301 25283 21335
rect 25225 21295 25283 21301
rect 25774 21292 25780 21344
rect 25832 21332 25838 21344
rect 25961 21335 26019 21341
rect 25961 21332 25973 21335
rect 25832 21304 25973 21332
rect 25832 21292 25838 21304
rect 25961 21301 25973 21304
rect 26007 21301 26019 21335
rect 25961 21295 26019 21301
rect 1104 21242 28152 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 28152 21242
rect 1104 21168 28152 21190
rect 3786 21088 3792 21140
rect 3844 21128 3850 21140
rect 3881 21131 3939 21137
rect 3881 21128 3893 21131
rect 3844 21100 3893 21128
rect 3844 21088 3850 21100
rect 3881 21097 3893 21100
rect 3927 21097 3939 21131
rect 3881 21091 3939 21097
rect 12342 21088 12348 21140
rect 12400 21088 12406 21140
rect 12710 21088 12716 21140
rect 12768 21128 12774 21140
rect 12805 21131 12863 21137
rect 12805 21128 12817 21131
rect 12768 21100 12817 21128
rect 12768 21088 12774 21100
rect 12805 21097 12817 21100
rect 12851 21128 12863 21131
rect 13998 21128 14004 21140
rect 12851 21100 14004 21128
rect 12851 21097 12863 21100
rect 12805 21091 12863 21097
rect 13998 21088 14004 21100
rect 14056 21088 14062 21140
rect 16298 21088 16304 21140
rect 16356 21128 16362 21140
rect 16485 21131 16543 21137
rect 16485 21128 16497 21131
rect 16356 21100 16497 21128
rect 16356 21088 16362 21100
rect 16485 21097 16497 21100
rect 16531 21097 16543 21131
rect 16485 21091 16543 21097
rect 17129 21131 17187 21137
rect 17129 21097 17141 21131
rect 17175 21128 17187 21131
rect 19058 21128 19064 21140
rect 17175 21100 19064 21128
rect 17175 21097 17187 21100
rect 17129 21091 17187 21097
rect 19058 21088 19064 21100
rect 19116 21088 19122 21140
rect 21174 21128 21180 21140
rect 19306 21100 21180 21128
rect 12728 21032 14872 21060
rect 6362 20952 6368 21004
rect 6420 20992 6426 21004
rect 6825 20995 6883 21001
rect 6420 20964 6684 20992
rect 6420 20952 6426 20964
rect 1026 20884 1032 20936
rect 1084 20924 1090 20936
rect 1949 20927 2007 20933
rect 1949 20924 1961 20927
rect 1084 20896 1961 20924
rect 1084 20884 1090 20896
rect 1949 20893 1961 20896
rect 1995 20893 2007 20927
rect 1949 20887 2007 20893
rect 2682 20884 2688 20936
rect 2740 20924 2746 20936
rect 3694 20924 3700 20936
rect 2740 20896 3700 20924
rect 2740 20884 2746 20896
rect 3694 20884 3700 20896
rect 3752 20924 3758 20936
rect 3789 20927 3847 20933
rect 3789 20924 3801 20927
rect 3752 20896 3801 20924
rect 3752 20884 3758 20896
rect 3789 20893 3801 20896
rect 3835 20893 3847 20927
rect 3789 20887 3847 20893
rect 3973 20927 4031 20933
rect 3973 20893 3985 20927
rect 4019 20924 4031 20927
rect 4062 20924 4068 20936
rect 4019 20896 4068 20924
rect 4019 20893 4031 20896
rect 3973 20887 4031 20893
rect 1486 20816 1492 20868
rect 1544 20816 1550 20868
rect 1762 20816 1768 20868
rect 1820 20856 1826 20868
rect 1857 20859 1915 20865
rect 1857 20856 1869 20859
rect 1820 20828 1869 20856
rect 1820 20816 1826 20828
rect 1857 20825 1869 20828
rect 1903 20856 1915 20859
rect 2130 20856 2136 20868
rect 1903 20828 2136 20856
rect 1903 20825 1915 20828
rect 1857 20819 1915 20825
rect 2130 20816 2136 20828
rect 2188 20816 2194 20868
rect 2225 20859 2283 20865
rect 2225 20825 2237 20859
rect 2271 20856 2283 20859
rect 2498 20856 2504 20868
rect 2271 20828 2504 20856
rect 2271 20825 2283 20828
rect 2225 20819 2283 20825
rect 2498 20816 2504 20828
rect 2556 20856 2562 20868
rect 3418 20856 3424 20868
rect 2556 20828 3424 20856
rect 2556 20816 2562 20828
rect 3418 20816 3424 20828
rect 3476 20816 3482 20868
rect 3804 20856 3832 20887
rect 4062 20884 4068 20896
rect 4120 20884 4126 20936
rect 4614 20884 4620 20936
rect 4672 20924 4678 20936
rect 4801 20927 4859 20933
rect 4801 20924 4813 20927
rect 4672 20896 4813 20924
rect 4672 20884 4678 20896
rect 4801 20893 4813 20896
rect 4847 20893 4859 20927
rect 4801 20887 4859 20893
rect 4982 20884 4988 20936
rect 5040 20884 5046 20936
rect 5626 20884 5632 20936
rect 5684 20884 5690 20936
rect 5718 20884 5724 20936
rect 5776 20884 5782 20936
rect 5905 20927 5963 20933
rect 5905 20893 5917 20927
rect 5951 20924 5963 20927
rect 6457 20927 6515 20933
rect 6457 20924 6469 20927
rect 5951 20896 6469 20924
rect 5951 20893 5963 20896
rect 5905 20887 5963 20893
rect 6457 20893 6469 20896
rect 6503 20893 6515 20927
rect 6656 20924 6684 20964
rect 6825 20961 6837 20995
rect 6871 20992 6883 20995
rect 7742 20992 7748 21004
rect 6871 20964 7748 20992
rect 6871 20961 6883 20964
rect 6825 20955 6883 20961
rect 7742 20952 7748 20964
rect 7800 20952 7806 21004
rect 6917 20927 6975 20933
rect 6917 20924 6929 20927
rect 6656 20896 6929 20924
rect 6457 20887 6515 20893
rect 6917 20893 6929 20896
rect 6963 20893 6975 20927
rect 6917 20887 6975 20893
rect 7101 20927 7159 20933
rect 7101 20893 7113 20927
rect 7147 20893 7159 20927
rect 7101 20887 7159 20893
rect 6472 20856 6500 20887
rect 7116 20856 7144 20887
rect 10594 20884 10600 20936
rect 10652 20884 10658 20936
rect 12728 20933 12756 21032
rect 12986 20952 12992 21004
rect 13044 20952 13050 21004
rect 12713 20927 12771 20933
rect 12713 20893 12725 20927
rect 12759 20893 12771 20927
rect 12713 20887 12771 20893
rect 13078 20884 13084 20936
rect 13136 20884 13142 20936
rect 13173 20927 13231 20933
rect 13173 20893 13185 20927
rect 13219 20893 13231 20927
rect 13173 20887 13231 20893
rect 13265 20927 13323 20933
rect 13265 20893 13277 20927
rect 13311 20924 13323 20927
rect 14093 20927 14151 20933
rect 14093 20924 14105 20927
rect 13311 20896 14105 20924
rect 13311 20893 13323 20896
rect 13265 20887 13323 20893
rect 14093 20893 14105 20896
rect 14139 20893 14151 20927
rect 14093 20887 14151 20893
rect 3804 20828 4108 20856
rect 6472 20828 7144 20856
rect 10873 20859 10931 20865
rect 4080 20800 4108 20828
rect 10873 20825 10885 20859
rect 10919 20856 10931 20859
rect 11146 20856 11152 20868
rect 10919 20828 11152 20856
rect 10919 20825 10931 20828
rect 10873 20819 10931 20825
rect 11146 20816 11152 20828
rect 11204 20816 11210 20868
rect 12250 20856 12256 20868
rect 12098 20828 12256 20856
rect 12250 20816 12256 20828
rect 12308 20816 12314 20868
rect 12986 20816 12992 20868
rect 13044 20856 13050 20868
rect 13188 20856 13216 20887
rect 14182 20884 14188 20936
rect 14240 20924 14246 20936
rect 14277 20927 14335 20933
rect 14277 20924 14289 20927
rect 14240 20896 14289 20924
rect 14240 20884 14246 20896
rect 14277 20893 14289 20896
rect 14323 20893 14335 20927
rect 14277 20887 14335 20893
rect 14366 20884 14372 20936
rect 14424 20924 14430 20936
rect 14461 20927 14519 20933
rect 14461 20924 14473 20927
rect 14424 20896 14473 20924
rect 14424 20884 14430 20896
rect 14461 20893 14473 20896
rect 14507 20893 14519 20927
rect 14461 20887 14519 20893
rect 14553 20927 14611 20933
rect 14553 20893 14565 20927
rect 14599 20924 14611 20927
rect 14642 20924 14648 20936
rect 14599 20896 14648 20924
rect 14599 20893 14611 20896
rect 14553 20887 14611 20893
rect 14642 20884 14648 20896
rect 14700 20884 14706 20936
rect 13044 20828 13216 20856
rect 13817 20859 13875 20865
rect 13044 20816 13050 20828
rect 13817 20825 13829 20859
rect 13863 20856 13875 20859
rect 14844 20856 14872 21032
rect 15102 21020 15108 21072
rect 15160 21060 15166 21072
rect 17862 21060 17868 21072
rect 15160 21032 15332 21060
rect 15160 21020 15166 21032
rect 15194 20952 15200 21004
rect 15252 20952 15258 21004
rect 15102 20884 15108 20936
rect 15160 20884 15166 20936
rect 15304 20924 15332 21032
rect 17696 21032 17868 21060
rect 16206 20952 16212 21004
rect 16264 20992 16270 21004
rect 16669 20995 16727 21001
rect 16669 20992 16681 20995
rect 16264 20964 16681 20992
rect 16264 20952 16270 20964
rect 16669 20961 16681 20964
rect 16715 20961 16727 20995
rect 16669 20955 16727 20961
rect 17126 20952 17132 21004
rect 17184 20992 17190 21004
rect 17313 20995 17371 21001
rect 17313 20992 17325 20995
rect 17184 20964 17325 20992
rect 17184 20952 17190 20964
rect 17313 20961 17325 20964
rect 17359 20961 17371 20995
rect 17313 20955 17371 20961
rect 17402 20952 17408 21004
rect 17460 20952 17466 21004
rect 17696 21001 17724 21032
rect 17862 21020 17868 21032
rect 17920 21020 17926 21072
rect 18598 21020 18604 21072
rect 18656 21060 18662 21072
rect 19306 21060 19334 21100
rect 21174 21088 21180 21100
rect 21232 21088 21238 21140
rect 23569 21131 23627 21137
rect 21652 21100 23244 21128
rect 18656 21032 19334 21060
rect 18656 21020 18662 21032
rect 19518 21020 19524 21072
rect 19576 21020 19582 21072
rect 19610 21020 19616 21072
rect 19668 21020 19674 21072
rect 21358 21060 21364 21072
rect 20916 21032 21364 21060
rect 17681 20995 17739 21001
rect 17681 20961 17693 20995
rect 17727 20961 17739 20995
rect 17681 20955 17739 20961
rect 17770 20952 17776 21004
rect 17828 20952 17834 21004
rect 17954 20952 17960 21004
rect 18012 20992 18018 21004
rect 20916 20992 20944 21032
rect 21358 21020 21364 21032
rect 21416 21020 21422 21072
rect 18012 20964 20944 20992
rect 21008 20964 21496 20992
rect 18012 20952 18018 20964
rect 15657 20927 15715 20933
rect 15657 20924 15669 20927
rect 15304 20896 15669 20924
rect 15657 20893 15669 20896
rect 15703 20893 15715 20927
rect 15657 20887 15715 20893
rect 16114 20884 16120 20936
rect 16172 20924 16178 20936
rect 16393 20927 16451 20933
rect 16393 20924 16405 20927
rect 16172 20896 16405 20924
rect 16172 20884 16178 20896
rect 16393 20893 16405 20896
rect 16439 20893 16451 20927
rect 16393 20887 16451 20893
rect 16574 20884 16580 20936
rect 16632 20924 16638 20936
rect 18598 20926 18604 20936
rect 18524 20924 18604 20926
rect 16632 20898 18604 20924
rect 16632 20896 18552 20898
rect 16632 20884 16638 20896
rect 18598 20884 18604 20898
rect 18656 20884 18662 20936
rect 18892 20933 18920 20964
rect 18877 20927 18935 20933
rect 18877 20893 18889 20927
rect 18923 20893 18935 20927
rect 18877 20887 18935 20893
rect 19058 20884 19064 20936
rect 19116 20924 19122 20936
rect 19245 20927 19303 20933
rect 19245 20924 19257 20927
rect 19116 20896 19257 20924
rect 19116 20884 19122 20896
rect 19245 20893 19257 20896
rect 19291 20893 19303 20927
rect 19245 20887 19303 20893
rect 19441 20927 19499 20933
rect 19441 20893 19453 20927
rect 19487 20924 19499 20927
rect 19610 20924 19616 20936
rect 19487 20896 19616 20924
rect 19487 20893 19499 20896
rect 19441 20887 19499 20893
rect 19610 20884 19616 20896
rect 19668 20884 19674 20936
rect 19705 20927 19763 20933
rect 19705 20893 19717 20927
rect 19751 20893 19763 20927
rect 19705 20887 19763 20893
rect 15470 20856 15476 20868
rect 13863 20828 14780 20856
rect 14844 20828 15476 20856
rect 13863 20825 13875 20828
rect 13817 20819 13875 20825
rect 4062 20748 4068 20800
rect 4120 20748 4126 20800
rect 4893 20791 4951 20797
rect 4893 20757 4905 20791
rect 4939 20788 4951 20791
rect 5261 20791 5319 20797
rect 5261 20788 5273 20791
rect 4939 20760 5273 20788
rect 4939 20757 4951 20760
rect 4893 20751 4951 20757
rect 5261 20757 5273 20760
rect 5307 20757 5319 20791
rect 5261 20751 5319 20757
rect 7098 20748 7104 20800
rect 7156 20748 7162 20800
rect 12526 20748 12532 20800
rect 12584 20748 12590 20800
rect 12618 20748 12624 20800
rect 12676 20788 12682 20800
rect 13354 20788 13360 20800
rect 12676 20760 13360 20788
rect 12676 20748 12682 20760
rect 13354 20748 13360 20760
rect 13412 20788 13418 20800
rect 13725 20791 13783 20797
rect 13725 20788 13737 20791
rect 13412 20760 13737 20788
rect 13412 20748 13418 20760
rect 13725 20757 13737 20760
rect 13771 20788 13783 20791
rect 13906 20788 13912 20800
rect 13771 20760 13912 20788
rect 13771 20757 13783 20760
rect 13725 20751 13783 20757
rect 13906 20748 13912 20760
rect 13964 20748 13970 20800
rect 14752 20788 14780 20828
rect 15470 20816 15476 20828
rect 15528 20816 15534 20868
rect 18322 20856 18328 20868
rect 16960 20828 18328 20856
rect 15838 20788 15844 20800
rect 14752 20760 15844 20788
rect 15838 20748 15844 20760
rect 15896 20748 15902 20800
rect 16960 20797 16988 20828
rect 18322 20816 18328 20828
rect 18380 20816 18386 20868
rect 18506 20816 18512 20868
rect 18564 20856 18570 20868
rect 18785 20859 18843 20865
rect 18785 20856 18797 20859
rect 18564 20828 18797 20856
rect 18564 20816 18570 20828
rect 18785 20825 18797 20828
rect 18831 20856 18843 20859
rect 19150 20856 19156 20868
rect 18831 20828 19156 20856
rect 18831 20825 18843 20828
rect 18785 20819 18843 20825
rect 19150 20816 19156 20828
rect 19208 20816 19214 20868
rect 19720 20856 19748 20887
rect 20070 20884 20076 20936
rect 20128 20884 20134 20936
rect 20162 20884 20168 20936
rect 20220 20884 20226 20936
rect 20530 20884 20536 20936
rect 20588 20924 20594 20936
rect 21008 20933 21036 20964
rect 20809 20927 20867 20933
rect 20809 20924 20821 20927
rect 20588 20896 20821 20924
rect 20588 20884 20594 20896
rect 20809 20893 20821 20896
rect 20855 20893 20867 20927
rect 20809 20887 20867 20893
rect 20993 20927 21051 20933
rect 20993 20893 21005 20927
rect 21039 20893 21051 20927
rect 20993 20887 21051 20893
rect 21082 20884 21088 20936
rect 21140 20924 21146 20936
rect 21468 20933 21496 20964
rect 21542 20952 21548 21004
rect 21600 20952 21606 21004
rect 21269 20927 21327 20933
rect 21269 20924 21281 20927
rect 21140 20896 21281 20924
rect 21140 20884 21146 20896
rect 21269 20893 21281 20896
rect 21315 20893 21327 20927
rect 21269 20887 21327 20893
rect 21453 20927 21511 20933
rect 21453 20893 21465 20927
rect 21499 20924 21511 20927
rect 21652 20924 21680 21100
rect 22002 21020 22008 21072
rect 22060 21060 22066 21072
rect 23109 21063 23167 21069
rect 23109 21060 23121 21063
rect 22060 21032 23121 21060
rect 22060 21020 22066 21032
rect 23109 21029 23121 21032
rect 23155 21029 23167 21063
rect 23216 21060 23244 21100
rect 23569 21097 23581 21131
rect 23615 21128 23627 21131
rect 23934 21128 23940 21140
rect 23615 21100 23940 21128
rect 23615 21097 23627 21100
rect 23569 21091 23627 21097
rect 23934 21088 23940 21100
rect 23992 21088 23998 21140
rect 25038 21088 25044 21140
rect 25096 21088 25102 21140
rect 26050 21088 26056 21140
rect 26108 21128 26114 21140
rect 27065 21131 27123 21137
rect 27065 21128 27077 21131
rect 26108 21100 27077 21128
rect 26108 21088 26114 21100
rect 27065 21097 27077 21100
rect 27111 21097 27123 21131
rect 27065 21091 27123 21097
rect 23216 21032 23428 21060
rect 23109 21023 23167 21029
rect 21729 20995 21787 21001
rect 21729 20961 21741 20995
rect 21775 20992 21787 20995
rect 22554 20992 22560 21004
rect 21775 20964 22560 20992
rect 21775 20961 21787 20964
rect 21729 20955 21787 20961
rect 22554 20952 22560 20964
rect 22612 20952 22618 21004
rect 23400 20936 23428 21032
rect 25056 20992 25084 21088
rect 25593 20995 25651 21001
rect 25593 20992 25605 20995
rect 25056 20964 25605 20992
rect 25593 20961 25605 20964
rect 25639 20961 25651 20995
rect 25593 20955 25651 20961
rect 21499 20896 21680 20924
rect 21821 20927 21879 20933
rect 21499 20893 21511 20896
rect 21453 20887 21511 20893
rect 21821 20893 21833 20927
rect 21867 20893 21879 20927
rect 21821 20887 21879 20893
rect 20254 20856 20260 20868
rect 19720 20828 20260 20856
rect 20254 20816 20260 20828
rect 20312 20816 20318 20868
rect 20717 20859 20775 20865
rect 20717 20825 20729 20859
rect 20763 20856 20775 20859
rect 21361 20859 21419 20865
rect 21361 20856 21373 20859
rect 20763 20828 21373 20856
rect 20763 20825 20775 20828
rect 20717 20819 20775 20825
rect 21361 20825 21373 20828
rect 21407 20825 21419 20859
rect 21836 20856 21864 20887
rect 22094 20884 22100 20936
rect 22152 20884 22158 20936
rect 22186 20884 22192 20936
rect 22244 20884 22250 20936
rect 22370 20884 22376 20936
rect 22428 20884 22434 20936
rect 22465 20927 22523 20933
rect 22465 20893 22477 20927
rect 22511 20893 22523 20927
rect 22465 20887 22523 20893
rect 21836 20828 22140 20856
rect 21361 20819 21419 20825
rect 16945 20791 17003 20797
rect 16945 20757 16957 20791
rect 16991 20757 17003 20791
rect 16945 20751 17003 20757
rect 17589 20791 17647 20797
rect 17589 20757 17601 20791
rect 17635 20788 17647 20791
rect 18046 20788 18052 20800
rect 17635 20760 18052 20788
rect 17635 20757 17647 20760
rect 17589 20751 17647 20757
rect 18046 20748 18052 20760
rect 18104 20748 18110 20800
rect 18417 20791 18475 20797
rect 18417 20757 18429 20791
rect 18463 20788 18475 20791
rect 18690 20788 18696 20800
rect 18463 20760 18696 20788
rect 18463 20757 18475 20760
rect 18417 20751 18475 20757
rect 18690 20748 18696 20760
rect 18748 20748 18754 20800
rect 19518 20748 19524 20800
rect 19576 20788 19582 20800
rect 19889 20791 19947 20797
rect 19889 20788 19901 20791
rect 19576 20760 19901 20788
rect 19576 20748 19582 20760
rect 19889 20757 19901 20760
rect 19935 20757 19947 20791
rect 19889 20751 19947 20757
rect 20346 20748 20352 20800
rect 20404 20748 20410 20800
rect 20898 20748 20904 20800
rect 20956 20788 20962 20800
rect 21545 20791 21603 20797
rect 21545 20788 21557 20791
rect 20956 20760 21557 20788
rect 20956 20748 20962 20760
rect 21545 20757 21557 20760
rect 21591 20757 21603 20791
rect 21545 20751 21603 20757
rect 21910 20748 21916 20800
rect 21968 20748 21974 20800
rect 22112 20788 22140 20828
rect 22278 20816 22284 20868
rect 22336 20856 22342 20868
rect 22480 20856 22508 20887
rect 22738 20884 22744 20936
rect 22796 20884 22802 20936
rect 23014 20884 23020 20936
rect 23072 20884 23078 20936
rect 23290 20884 23296 20936
rect 23348 20884 23354 20936
rect 23382 20884 23388 20936
rect 23440 20884 23446 20936
rect 24302 20924 24308 20936
rect 23485 20896 24308 20924
rect 23308 20856 23336 20884
rect 23485 20856 23513 20896
rect 24302 20884 24308 20896
rect 24360 20884 24366 20936
rect 24394 20884 24400 20936
rect 24452 20924 24458 20936
rect 25314 20924 25320 20936
rect 24452 20896 25320 20924
rect 24452 20884 24458 20896
rect 25314 20884 25320 20896
rect 25372 20884 25378 20936
rect 22336 20828 22968 20856
rect 23308 20828 23513 20856
rect 22336 20816 22342 20828
rect 22186 20788 22192 20800
rect 22112 20760 22192 20788
rect 22186 20748 22192 20760
rect 22244 20748 22250 20800
rect 22370 20748 22376 20800
rect 22428 20788 22434 20800
rect 22738 20788 22744 20800
rect 22428 20760 22744 20788
rect 22428 20748 22434 20760
rect 22738 20748 22744 20760
rect 22796 20748 22802 20800
rect 22940 20797 22968 20828
rect 23566 20816 23572 20868
rect 23624 20816 23630 20868
rect 24857 20859 24915 20865
rect 24857 20825 24869 20859
rect 24903 20856 24915 20859
rect 25866 20856 25872 20868
rect 24903 20828 25872 20856
rect 24903 20825 24915 20828
rect 24857 20819 24915 20825
rect 25866 20816 25872 20828
rect 25924 20816 25930 20868
rect 26602 20816 26608 20868
rect 26660 20816 26666 20868
rect 22925 20791 22983 20797
rect 22925 20757 22937 20791
rect 22971 20788 22983 20791
rect 24210 20788 24216 20800
rect 22971 20760 24216 20788
rect 22971 20757 22983 20760
rect 22925 20751 22983 20757
rect 24210 20748 24216 20760
rect 24268 20748 24274 20800
rect 25038 20748 25044 20800
rect 25096 20797 25102 20800
rect 25096 20791 25115 20797
rect 25103 20757 25115 20791
rect 25096 20751 25115 20757
rect 25096 20748 25102 20751
rect 25222 20748 25228 20800
rect 25280 20748 25286 20800
rect 1104 20698 28152 20720
rect 1104 20646 4874 20698
rect 4926 20646 4938 20698
rect 4990 20646 5002 20698
rect 5054 20646 5066 20698
rect 5118 20646 5130 20698
rect 5182 20646 28152 20698
rect 1104 20624 28152 20646
rect 7653 20587 7711 20593
rect 7653 20553 7665 20587
rect 7699 20584 7711 20587
rect 8386 20584 8392 20596
rect 7699 20556 8392 20584
rect 7699 20553 7711 20556
rect 7653 20547 7711 20553
rect 8386 20544 8392 20556
rect 8444 20544 8450 20596
rect 11146 20544 11152 20596
rect 11204 20584 11210 20596
rect 11609 20587 11667 20593
rect 11609 20584 11621 20587
rect 11204 20556 11621 20584
rect 11204 20544 11210 20556
rect 11609 20553 11621 20556
rect 11655 20553 11667 20587
rect 12710 20584 12716 20596
rect 11609 20547 11667 20553
rect 12176 20556 12716 20584
rect 1946 20476 1952 20528
rect 2004 20476 2010 20528
rect 4154 20476 4160 20528
rect 4212 20516 4218 20528
rect 4212 20488 5028 20516
rect 4212 20476 4218 20488
rect 2596 20460 2648 20466
rect 2682 20408 2688 20460
rect 2740 20408 2746 20460
rect 4798 20408 4804 20460
rect 4856 20408 4862 20460
rect 5000 20457 5028 20488
rect 7098 20476 7104 20528
rect 7156 20476 7162 20528
rect 4985 20451 5043 20457
rect 4985 20417 4997 20451
rect 5031 20417 5043 20451
rect 4985 20411 5043 20417
rect 5718 20408 5724 20460
rect 5776 20408 5782 20460
rect 7558 20408 7564 20460
rect 7616 20448 7622 20460
rect 7653 20451 7711 20457
rect 7653 20448 7665 20451
rect 7616 20420 7665 20448
rect 7616 20408 7622 20420
rect 7653 20417 7665 20420
rect 7699 20417 7711 20451
rect 7653 20411 7711 20417
rect 11701 20451 11759 20457
rect 11701 20417 11713 20451
rect 11747 20448 11759 20451
rect 12176 20448 12204 20556
rect 12710 20544 12716 20556
rect 12768 20544 12774 20596
rect 12989 20587 13047 20593
rect 12989 20553 13001 20587
rect 13035 20584 13047 20587
rect 13078 20584 13084 20596
rect 13035 20556 13084 20584
rect 13035 20553 13047 20556
rect 12989 20547 13047 20553
rect 13078 20544 13084 20556
rect 13136 20544 13142 20596
rect 14737 20587 14795 20593
rect 13280 20556 14044 20584
rect 12526 20476 12532 20528
rect 12584 20476 12590 20528
rect 13280 20516 13308 20556
rect 13188 20488 13308 20516
rect 13464 20488 13768 20516
rect 11747 20420 12204 20448
rect 12253 20451 12311 20457
rect 11747 20417 11759 20420
rect 11701 20411 11759 20417
rect 12253 20417 12265 20451
rect 12299 20448 12311 20451
rect 12544 20448 12572 20476
rect 12299 20420 12572 20448
rect 12621 20451 12679 20457
rect 12299 20417 12311 20420
rect 12253 20411 12311 20417
rect 12621 20417 12633 20451
rect 12667 20417 12679 20451
rect 12621 20411 12679 20417
rect 2596 20402 2648 20408
rect 4893 20383 4951 20389
rect 4893 20349 4905 20383
rect 4939 20380 4951 20383
rect 5353 20383 5411 20389
rect 5353 20380 5365 20383
rect 4939 20352 5365 20380
rect 4939 20349 4951 20352
rect 4893 20343 4951 20349
rect 5353 20349 5365 20352
rect 5399 20380 5411 20383
rect 5626 20380 5632 20392
rect 5399 20352 5632 20380
rect 5399 20349 5411 20352
rect 5353 20343 5411 20349
rect 5626 20340 5632 20352
rect 5684 20340 5690 20392
rect 6181 20383 6239 20389
rect 6181 20349 6193 20383
rect 6227 20380 6239 20383
rect 6454 20380 6460 20392
rect 6227 20352 6460 20380
rect 6227 20349 6239 20352
rect 6181 20343 6239 20349
rect 6454 20340 6460 20352
rect 6512 20340 6518 20392
rect 7742 20340 7748 20392
rect 7800 20340 7806 20392
rect 11790 20340 11796 20392
rect 11848 20340 11854 20392
rect 12342 20340 12348 20392
rect 12400 20340 12406 20392
rect 12529 20383 12587 20389
rect 12529 20349 12541 20383
rect 12575 20349 12587 20383
rect 12636 20380 12664 20411
rect 12710 20408 12716 20460
rect 12768 20448 12774 20460
rect 13188 20457 13216 20488
rect 13464 20460 13492 20488
rect 13173 20451 13231 20457
rect 13173 20448 13185 20451
rect 12768 20420 13185 20448
rect 12768 20408 12774 20420
rect 13173 20417 13185 20420
rect 13219 20417 13231 20451
rect 13173 20411 13231 20417
rect 13265 20451 13323 20457
rect 13265 20417 13277 20451
rect 13311 20448 13323 20451
rect 13354 20448 13360 20460
rect 13311 20420 13360 20448
rect 13311 20417 13323 20420
rect 13265 20411 13323 20417
rect 13354 20408 13360 20420
rect 13412 20408 13418 20460
rect 13446 20408 13452 20460
rect 13504 20408 13510 20460
rect 13538 20408 13544 20460
rect 13596 20408 13602 20460
rect 13740 20457 13768 20488
rect 13633 20451 13691 20457
rect 13633 20417 13645 20451
rect 13679 20417 13691 20451
rect 13633 20411 13691 20417
rect 13725 20451 13783 20457
rect 13725 20417 13737 20451
rect 13771 20417 13783 20451
rect 13725 20411 13783 20417
rect 12802 20380 12808 20392
rect 12636 20352 12808 20380
rect 12529 20343 12587 20349
rect 11885 20315 11943 20321
rect 11885 20281 11897 20315
rect 11931 20312 11943 20315
rect 11974 20312 11980 20324
rect 11931 20284 11980 20312
rect 11931 20281 11943 20284
rect 11885 20275 11943 20281
rect 11974 20272 11980 20284
rect 12032 20272 12038 20324
rect 12434 20272 12440 20324
rect 12492 20312 12498 20324
rect 12544 20312 12572 20343
rect 12802 20340 12808 20352
rect 12860 20380 12866 20392
rect 13648 20380 13676 20411
rect 13906 20408 13912 20460
rect 13964 20408 13970 20460
rect 14016 20457 14044 20556
rect 14737 20553 14749 20587
rect 14783 20584 14795 20587
rect 15010 20584 15016 20596
rect 14783 20556 15016 20584
rect 14783 20553 14795 20556
rect 14737 20547 14795 20553
rect 15010 20544 15016 20556
rect 15068 20544 15074 20596
rect 15562 20544 15568 20596
rect 15620 20584 15626 20596
rect 16025 20587 16083 20593
rect 16025 20584 16037 20587
rect 15620 20556 16037 20584
rect 15620 20544 15626 20556
rect 16025 20553 16037 20556
rect 16071 20553 16083 20587
rect 16025 20547 16083 20553
rect 16390 20544 16396 20596
rect 16448 20544 16454 20596
rect 19610 20584 19616 20596
rect 17604 20556 19616 20584
rect 14090 20476 14096 20528
rect 14148 20516 14154 20528
rect 14185 20519 14243 20525
rect 14185 20516 14197 20519
rect 14148 20488 14197 20516
rect 14148 20476 14154 20488
rect 14185 20485 14197 20488
rect 14231 20485 14243 20519
rect 14185 20479 14243 20485
rect 15933 20519 15991 20525
rect 15933 20485 15945 20519
rect 15979 20516 15991 20519
rect 16298 20516 16304 20528
rect 15979 20488 16304 20516
rect 15979 20485 15991 20488
rect 15933 20479 15991 20485
rect 16298 20476 16304 20488
rect 16356 20476 16362 20528
rect 16408 20516 16436 20544
rect 16408 20488 16712 20516
rect 14001 20451 14059 20457
rect 14001 20417 14013 20451
rect 14047 20417 14059 20451
rect 14001 20411 14059 20417
rect 12860 20352 13216 20380
rect 12860 20340 12866 20352
rect 13078 20312 13084 20324
rect 12492 20284 13084 20312
rect 12492 20272 12498 20284
rect 13078 20272 13084 20284
rect 13136 20272 13142 20324
rect 13188 20312 13216 20352
rect 13556 20352 13676 20380
rect 13556 20312 13584 20352
rect 13188 20284 13584 20312
rect 14016 20312 14044 20411
rect 14550 20408 14556 20460
rect 14608 20408 14614 20460
rect 15286 20408 15292 20460
rect 15344 20408 15350 20460
rect 15378 20408 15384 20460
rect 15436 20408 15442 20460
rect 16206 20408 16212 20460
rect 16264 20408 16270 20460
rect 16684 20457 16712 20488
rect 16669 20451 16727 20457
rect 16669 20417 16681 20451
rect 16715 20417 16727 20451
rect 16669 20411 16727 20417
rect 17034 20408 17040 20460
rect 17092 20408 17098 20460
rect 17604 20457 17632 20556
rect 19610 20544 19616 20556
rect 19668 20544 19674 20596
rect 19886 20544 19892 20596
rect 19944 20584 19950 20596
rect 20993 20587 21051 20593
rect 19944 20556 20852 20584
rect 19944 20544 19950 20556
rect 18506 20516 18512 20528
rect 18340 20488 18512 20516
rect 17589 20451 17647 20457
rect 17589 20417 17601 20451
rect 17635 20417 17647 20451
rect 17589 20411 17647 20417
rect 17678 20408 17684 20460
rect 17736 20408 17742 20460
rect 18340 20457 18368 20488
rect 18506 20476 18512 20488
rect 18564 20476 18570 20528
rect 19518 20476 19524 20528
rect 19576 20476 19582 20528
rect 20824 20516 20852 20556
rect 20993 20553 21005 20587
rect 21039 20584 21051 20587
rect 21082 20584 21088 20596
rect 21039 20556 21088 20584
rect 21039 20553 21051 20556
rect 20993 20547 21051 20553
rect 21082 20544 21088 20556
rect 21140 20544 21146 20596
rect 22002 20544 22008 20596
rect 22060 20593 22066 20596
rect 22060 20587 22079 20593
rect 22067 20553 22079 20587
rect 22060 20547 22079 20553
rect 22060 20544 22066 20547
rect 22186 20544 22192 20596
rect 22244 20544 22250 20596
rect 24210 20544 24216 20596
rect 24268 20544 24274 20596
rect 25038 20544 25044 20596
rect 25096 20584 25102 20596
rect 25593 20587 25651 20593
rect 25593 20584 25605 20587
rect 25096 20556 25605 20584
rect 25096 20544 25102 20556
rect 25593 20553 25605 20556
rect 25639 20584 25651 20587
rect 25866 20584 25872 20596
rect 25639 20556 25872 20584
rect 25639 20553 25651 20556
rect 25593 20547 25651 20553
rect 25866 20544 25872 20556
rect 25924 20544 25930 20596
rect 26234 20544 26240 20596
rect 26292 20584 26298 20596
rect 26421 20587 26479 20593
rect 26421 20584 26433 20587
rect 26292 20556 26433 20584
rect 26292 20544 26298 20556
rect 26421 20553 26433 20556
rect 26467 20553 26479 20587
rect 26421 20547 26479 20553
rect 21269 20519 21327 20525
rect 21269 20516 21281 20519
rect 20824 20488 21281 20516
rect 21269 20485 21281 20488
rect 21315 20485 21327 20519
rect 21269 20479 21327 20485
rect 21818 20476 21824 20528
rect 21876 20476 21882 20528
rect 22830 20516 22836 20528
rect 22296 20488 22836 20516
rect 18325 20451 18383 20457
rect 18325 20417 18337 20451
rect 18371 20417 18383 20451
rect 18325 20411 18383 20417
rect 18785 20451 18843 20457
rect 18785 20417 18797 20451
rect 18831 20417 18843 20451
rect 18785 20411 18843 20417
rect 18877 20451 18935 20457
rect 18877 20417 18889 20451
rect 18923 20417 18935 20451
rect 18877 20411 18935 20417
rect 19061 20451 19119 20457
rect 19061 20417 19073 20451
rect 19107 20417 19119 20451
rect 19061 20411 19119 20417
rect 14366 20340 14372 20392
rect 14424 20340 14430 20392
rect 16393 20383 16451 20389
rect 16393 20349 16405 20383
rect 16439 20380 16451 20383
rect 16439 20352 17080 20380
rect 16439 20349 16451 20352
rect 16393 20343 16451 20349
rect 17052 20321 17080 20352
rect 18230 20340 18236 20392
rect 18288 20380 18294 20392
rect 18800 20380 18828 20411
rect 18288 20352 18828 20380
rect 18892 20380 18920 20411
rect 19076 20380 19104 20411
rect 19150 20408 19156 20460
rect 19208 20408 19214 20460
rect 20622 20408 20628 20460
rect 20680 20408 20686 20460
rect 21085 20451 21143 20457
rect 21085 20417 21097 20451
rect 21131 20448 21143 20451
rect 21174 20448 21180 20460
rect 21131 20420 21180 20448
rect 21131 20417 21143 20420
rect 21085 20411 21143 20417
rect 21174 20408 21180 20420
rect 21232 20408 21238 20460
rect 21358 20408 21364 20460
rect 21416 20408 21422 20460
rect 22296 20457 22324 20488
rect 22830 20476 22836 20488
rect 22888 20476 22894 20528
rect 26513 20519 26571 20525
rect 26513 20485 26525 20519
rect 26559 20516 26571 20519
rect 26970 20516 26976 20528
rect 26559 20488 26976 20516
rect 26559 20485 26571 20488
rect 26513 20479 26571 20485
rect 26970 20476 26976 20488
rect 27028 20476 27034 20528
rect 22281 20451 22339 20457
rect 22281 20417 22293 20451
rect 22327 20417 22339 20451
rect 24121 20451 24179 20457
rect 24121 20448 24133 20451
rect 22281 20411 22339 20417
rect 18892 20352 18946 20380
rect 19076 20352 19196 20380
rect 18288 20340 18294 20352
rect 17037 20315 17095 20321
rect 14016 20284 15608 20312
rect 12802 20204 12808 20256
rect 12860 20244 12866 20256
rect 13446 20244 13452 20256
rect 12860 20216 13452 20244
rect 12860 20204 12866 20216
rect 13446 20204 13452 20216
rect 13504 20204 13510 20256
rect 15580 20244 15608 20284
rect 17037 20281 17049 20315
rect 17083 20312 17095 20315
rect 17126 20312 17132 20324
rect 17083 20284 17132 20312
rect 17083 20281 17095 20284
rect 17037 20275 17095 20281
rect 17126 20272 17132 20284
rect 17184 20272 17190 20324
rect 17310 20272 17316 20324
rect 17368 20312 17374 20324
rect 17368 20284 18736 20312
rect 17368 20272 17374 20284
rect 18230 20244 18236 20256
rect 15580 20216 18236 20244
rect 18230 20204 18236 20216
rect 18288 20204 18294 20256
rect 18506 20204 18512 20256
rect 18564 20244 18570 20256
rect 18601 20247 18659 20253
rect 18601 20244 18613 20247
rect 18564 20216 18613 20244
rect 18564 20204 18570 20216
rect 18601 20213 18613 20216
rect 18647 20213 18659 20247
rect 18708 20244 18736 20284
rect 18918 20244 18946 20352
rect 19168 20324 19196 20352
rect 19242 20340 19248 20392
rect 19300 20340 19306 20392
rect 22554 20340 22560 20392
rect 22612 20340 22618 20392
rect 19150 20272 19156 20324
rect 19208 20272 19214 20324
rect 20622 20272 20628 20324
rect 20680 20312 20686 20324
rect 20680 20284 22416 20312
rect 20680 20272 20686 20284
rect 19886 20244 19892 20256
rect 18708 20216 19892 20244
rect 18601 20207 18659 20213
rect 19886 20204 19892 20216
rect 19944 20204 19950 20256
rect 20070 20204 20076 20256
rect 20128 20244 20134 20256
rect 21085 20247 21143 20253
rect 21085 20244 21097 20247
rect 20128 20216 21097 20244
rect 20128 20204 20134 20216
rect 21085 20213 21097 20216
rect 21131 20213 21143 20247
rect 21085 20207 21143 20213
rect 21910 20204 21916 20256
rect 21968 20244 21974 20256
rect 22005 20247 22063 20253
rect 22005 20244 22017 20247
rect 21968 20216 22017 20244
rect 21968 20204 21974 20216
rect 22005 20213 22017 20216
rect 22051 20213 22063 20247
rect 22388 20244 22416 20284
rect 23676 20244 23704 20434
rect 24044 20420 24133 20448
rect 24044 20256 24072 20420
rect 24121 20417 24133 20420
rect 24167 20417 24179 20451
rect 24121 20411 24179 20417
rect 25774 20408 25780 20460
rect 25832 20408 25838 20460
rect 26053 20451 26111 20457
rect 26053 20417 26065 20451
rect 26099 20448 26111 20451
rect 26142 20448 26148 20460
rect 26099 20420 26148 20448
rect 26099 20417 26111 20420
rect 26053 20411 26111 20417
rect 26142 20408 26148 20420
rect 26200 20408 26206 20460
rect 26234 20408 26240 20460
rect 26292 20408 26298 20460
rect 23750 20244 23756 20256
rect 22388 20216 23756 20244
rect 22005 20207 22063 20213
rect 23750 20204 23756 20216
rect 23808 20204 23814 20256
rect 24026 20204 24032 20256
rect 24084 20204 24090 20256
rect 1104 20154 28152 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 28152 20154
rect 1104 20080 28152 20102
rect 4341 20043 4399 20049
rect 4341 20009 4353 20043
rect 4387 20040 4399 20043
rect 4798 20040 4804 20052
rect 4387 20012 4804 20040
rect 4387 20009 4399 20012
rect 4341 20003 4399 20009
rect 4798 20000 4804 20012
rect 4856 20000 4862 20052
rect 12342 20000 12348 20052
rect 12400 20040 12406 20052
rect 13081 20043 13139 20049
rect 13081 20040 13093 20043
rect 12400 20012 13093 20040
rect 12400 20000 12406 20012
rect 13081 20009 13093 20012
rect 13127 20009 13139 20043
rect 13081 20003 13139 20009
rect 14553 20043 14611 20049
rect 14553 20009 14565 20043
rect 14599 20040 14611 20043
rect 14918 20040 14924 20052
rect 14599 20012 14924 20040
rect 14599 20009 14611 20012
rect 14553 20003 14611 20009
rect 14918 20000 14924 20012
rect 14976 20000 14982 20052
rect 15194 20000 15200 20052
rect 15252 20000 15258 20052
rect 15470 20000 15476 20052
rect 15528 20000 15534 20052
rect 16206 20000 16212 20052
rect 16264 20040 16270 20052
rect 16577 20043 16635 20049
rect 16577 20040 16589 20043
rect 16264 20012 16589 20040
rect 16264 20000 16270 20012
rect 16577 20009 16589 20012
rect 16623 20009 16635 20043
rect 16577 20003 16635 20009
rect 18230 20000 18236 20052
rect 18288 20040 18294 20052
rect 22465 20043 22523 20049
rect 18288 20012 22140 20040
rect 18288 20000 18294 20012
rect 22112 19984 22140 20012
rect 22465 20009 22477 20043
rect 22511 20040 22523 20043
rect 22554 20040 22560 20052
rect 22511 20012 22560 20040
rect 22511 20009 22523 20012
rect 22465 20003 22523 20009
rect 22554 20000 22560 20012
rect 22612 20000 22618 20052
rect 23382 20000 23388 20052
rect 23440 20040 23446 20052
rect 23661 20043 23719 20049
rect 23661 20040 23673 20043
rect 23440 20012 23673 20040
rect 23440 20000 23446 20012
rect 23661 20009 23673 20012
rect 23707 20009 23719 20043
rect 23661 20003 23719 20009
rect 23845 20043 23903 20049
rect 23845 20009 23857 20043
rect 23891 20009 23903 20043
rect 23845 20003 23903 20009
rect 1578 19932 1584 19984
rect 1636 19972 1642 19984
rect 9122 19972 9128 19984
rect 1636 19944 9128 19972
rect 1636 19932 1642 19944
rect 9122 19932 9128 19944
rect 9180 19932 9186 19984
rect 12437 19975 12495 19981
rect 12437 19941 12449 19975
rect 12483 19972 12495 19975
rect 13262 19972 13268 19984
rect 12483 19944 13268 19972
rect 12483 19941 12495 19944
rect 12437 19935 12495 19941
rect 13262 19932 13268 19944
rect 13320 19932 13326 19984
rect 14642 19972 14648 19984
rect 13464 19944 14648 19972
rect 2133 19907 2191 19913
rect 2133 19873 2145 19907
rect 2179 19904 2191 19907
rect 7653 19907 7711 19913
rect 2179 19876 2452 19904
rect 2179 19873 2191 19876
rect 2133 19867 2191 19873
rect 2424 19848 2452 19876
rect 7653 19873 7665 19907
rect 7699 19904 7711 19907
rect 7742 19904 7748 19916
rect 7699 19876 7748 19904
rect 7699 19873 7711 19876
rect 7653 19867 7711 19873
rect 7742 19864 7748 19876
rect 7800 19864 7806 19916
rect 10594 19864 10600 19916
rect 10652 19904 10658 19916
rect 10689 19907 10747 19913
rect 10689 19904 10701 19907
rect 10652 19876 10701 19904
rect 10652 19864 10658 19876
rect 10689 19873 10701 19876
rect 10735 19873 10747 19907
rect 10689 19867 10747 19873
rect 10965 19907 11023 19913
rect 10965 19873 10977 19907
rect 11011 19904 11023 19907
rect 11974 19904 11980 19916
rect 11011 19876 11980 19904
rect 11011 19873 11023 19876
rect 10965 19867 11023 19873
rect 11974 19864 11980 19876
rect 12032 19864 12038 19916
rect 12529 19907 12587 19913
rect 12529 19873 12541 19907
rect 12575 19904 12587 19907
rect 12618 19904 12624 19916
rect 12575 19876 12624 19904
rect 12575 19873 12587 19876
rect 12529 19867 12587 19873
rect 12618 19864 12624 19876
rect 12676 19864 12682 19916
rect 12710 19864 12716 19916
rect 12768 19864 12774 19916
rect 12989 19907 13047 19913
rect 12989 19873 13001 19907
rect 13035 19904 13047 19907
rect 13078 19904 13084 19916
rect 13035 19876 13084 19904
rect 13035 19873 13047 19876
rect 12989 19867 13047 19873
rect 13078 19864 13084 19876
rect 13136 19904 13142 19916
rect 13464 19904 13492 19944
rect 14642 19932 14648 19944
rect 14700 19972 14706 19984
rect 19334 19972 19340 19984
rect 14700 19944 15332 19972
rect 14700 19932 14706 19944
rect 13136 19876 13492 19904
rect 13556 19876 13768 19904
rect 13136 19864 13142 19876
rect 842 19796 848 19848
rect 900 19836 906 19848
rect 1397 19839 1455 19845
rect 1397 19836 1409 19839
rect 900 19808 1409 19836
rect 900 19796 906 19808
rect 1397 19805 1409 19808
rect 1443 19805 1455 19839
rect 1397 19799 1455 19805
rect 1946 19796 1952 19848
rect 2004 19836 2010 19848
rect 2041 19839 2099 19845
rect 2041 19836 2053 19839
rect 2004 19808 2053 19836
rect 2004 19796 2010 19808
rect 2041 19805 2053 19808
rect 2087 19805 2099 19839
rect 2041 19799 2099 19805
rect 2222 19796 2228 19848
rect 2280 19796 2286 19848
rect 2406 19796 2412 19848
rect 2464 19796 2470 19848
rect 2866 19796 2872 19848
rect 2924 19796 2930 19848
rect 4154 19796 4160 19848
rect 4212 19836 4218 19848
rect 4249 19839 4307 19845
rect 4249 19836 4261 19839
rect 4212 19808 4261 19836
rect 4212 19796 4218 19808
rect 4249 19805 4261 19808
rect 4295 19836 4307 19839
rect 5350 19836 5356 19848
rect 4295 19808 5356 19836
rect 4295 19805 4307 19808
rect 4249 19799 4307 19805
rect 5350 19796 5356 19808
rect 5408 19836 5414 19848
rect 7374 19836 7380 19848
rect 5408 19808 7380 19836
rect 5408 19796 5414 19808
rect 7374 19796 7380 19808
rect 7432 19796 7438 19848
rect 7558 19796 7564 19848
rect 7616 19796 7622 19848
rect 8110 19796 8116 19848
rect 8168 19836 8174 19848
rect 9033 19839 9091 19845
rect 9033 19836 9045 19839
rect 8168 19808 9045 19836
rect 8168 19796 8174 19808
rect 9033 19805 9045 19808
rect 9079 19805 9091 19839
rect 9033 19799 9091 19805
rect 9217 19839 9275 19845
rect 9217 19805 9229 19839
rect 9263 19805 9275 19839
rect 9217 19799 9275 19805
rect 12897 19839 12955 19845
rect 12897 19805 12909 19839
rect 12943 19836 12955 19839
rect 13173 19839 13231 19845
rect 13173 19836 13185 19839
rect 12943 19808 13185 19836
rect 12943 19805 12955 19808
rect 12897 19799 12955 19805
rect 13173 19805 13185 19808
rect 13219 19805 13231 19839
rect 13173 19799 13231 19805
rect 1673 19771 1731 19777
rect 1673 19737 1685 19771
rect 1719 19768 1731 19771
rect 2682 19768 2688 19780
rect 1719 19740 2688 19768
rect 1719 19737 1731 19740
rect 1673 19731 1731 19737
rect 2682 19728 2688 19740
rect 2740 19728 2746 19780
rect 3421 19771 3479 19777
rect 3421 19737 3433 19771
rect 3467 19768 3479 19771
rect 3694 19768 3700 19780
rect 3467 19740 3700 19768
rect 3467 19737 3479 19740
rect 3421 19731 3479 19737
rect 3694 19728 3700 19740
rect 3752 19728 3758 19780
rect 8386 19728 8392 19780
rect 8444 19768 8450 19780
rect 9232 19768 9260 19799
rect 13262 19796 13268 19848
rect 13320 19836 13326 19848
rect 13357 19839 13415 19845
rect 13357 19836 13369 19839
rect 13320 19808 13369 19836
rect 13320 19796 13326 19808
rect 13357 19805 13369 19808
rect 13403 19805 13415 19839
rect 13357 19799 13415 19805
rect 12250 19768 12256 19780
rect 8444 19740 9260 19768
rect 12190 19740 12256 19768
rect 8444 19728 8450 19740
rect 12250 19728 12256 19740
rect 12308 19728 12314 19780
rect 12805 19771 12863 19777
rect 12805 19737 12817 19771
rect 12851 19737 12863 19771
rect 13372 19768 13400 19799
rect 13446 19796 13452 19848
rect 13504 19836 13510 19848
rect 13556 19845 13584 19876
rect 13740 19848 13768 19876
rect 15010 19864 15016 19916
rect 15068 19904 15074 19916
rect 15197 19907 15255 19913
rect 15197 19904 15209 19907
rect 15068 19876 15209 19904
rect 15068 19864 15074 19876
rect 15197 19873 15209 19876
rect 15243 19873 15255 19907
rect 15304 19904 15332 19944
rect 19260 19944 19340 19972
rect 17954 19904 17960 19916
rect 15304 19876 17960 19904
rect 15197 19867 15255 19873
rect 13541 19839 13599 19845
rect 13541 19836 13553 19839
rect 13504 19808 13553 19836
rect 13504 19796 13510 19808
rect 13541 19805 13553 19808
rect 13587 19805 13599 19839
rect 13541 19799 13599 19805
rect 13633 19839 13691 19845
rect 13633 19805 13645 19839
rect 13679 19805 13691 19839
rect 13633 19799 13691 19805
rect 13648 19768 13676 19799
rect 13722 19796 13728 19848
rect 13780 19836 13786 19848
rect 13817 19839 13875 19845
rect 13817 19836 13829 19839
rect 13780 19808 13829 19836
rect 13780 19796 13786 19808
rect 13817 19805 13829 19808
rect 13863 19805 13875 19839
rect 13817 19799 13875 19805
rect 13906 19796 13912 19848
rect 13964 19836 13970 19848
rect 14366 19836 14372 19848
rect 13964 19808 14372 19836
rect 13964 19796 13970 19808
rect 14366 19796 14372 19808
rect 14424 19796 14430 19848
rect 14550 19796 14556 19848
rect 14608 19796 14614 19848
rect 15102 19796 15108 19848
rect 15160 19796 15166 19848
rect 16316 19845 16344 19876
rect 17954 19864 17960 19876
rect 18012 19864 18018 19916
rect 18708 19876 18920 19904
rect 16301 19839 16359 19845
rect 16301 19805 16313 19839
rect 16347 19805 16359 19839
rect 16301 19799 16359 19805
rect 16390 19796 16396 19848
rect 16448 19796 16454 19848
rect 18708 19845 18736 19876
rect 18601 19839 18659 19845
rect 18601 19805 18613 19839
rect 18647 19805 18659 19839
rect 18601 19799 18659 19805
rect 18693 19839 18751 19845
rect 18693 19805 18705 19839
rect 18739 19805 18751 19839
rect 18693 19799 18751 19805
rect 16574 19768 16580 19780
rect 13372 19740 13676 19768
rect 16408 19740 16580 19768
rect 12805 19731 12863 19737
rect 7834 19660 7840 19712
rect 7892 19700 7898 19712
rect 7929 19703 7987 19709
rect 7929 19700 7941 19703
rect 7892 19672 7941 19700
rect 7892 19660 7898 19672
rect 7929 19669 7941 19672
rect 7975 19669 7987 19703
rect 7929 19663 7987 19669
rect 10042 19660 10048 19712
rect 10100 19660 10106 19712
rect 12820 19700 12848 19731
rect 16408 19712 16436 19740
rect 16574 19728 16580 19740
rect 16632 19728 16638 19780
rect 16758 19728 16764 19780
rect 16816 19768 16822 19780
rect 17218 19768 17224 19780
rect 16816 19740 17224 19768
rect 16816 19728 16822 19740
rect 17218 19728 17224 19740
rect 17276 19768 17282 19780
rect 17957 19771 18015 19777
rect 17957 19768 17969 19771
rect 17276 19740 17969 19768
rect 17276 19728 17282 19740
rect 17957 19737 17969 19740
rect 18003 19737 18015 19771
rect 17957 19731 18015 19737
rect 12894 19700 12900 19712
rect 12820 19672 12900 19700
rect 12894 19660 12900 19672
rect 12952 19700 12958 19712
rect 13633 19703 13691 19709
rect 13633 19700 13645 19703
rect 12952 19672 13645 19700
rect 12952 19660 12958 19672
rect 13633 19669 13645 19672
rect 13679 19669 13691 19703
rect 13633 19663 13691 19669
rect 16390 19660 16396 19712
rect 16448 19660 16454 19712
rect 18138 19660 18144 19712
rect 18196 19700 18202 19712
rect 18417 19703 18475 19709
rect 18417 19700 18429 19703
rect 18196 19672 18429 19700
rect 18196 19660 18202 19672
rect 18417 19669 18429 19672
rect 18463 19669 18475 19703
rect 18616 19700 18644 19799
rect 18782 19796 18788 19848
rect 18840 19796 18846 19848
rect 18892 19836 18920 19876
rect 18966 19864 18972 19916
rect 19024 19904 19030 19916
rect 19061 19907 19119 19913
rect 19061 19904 19073 19907
rect 19024 19876 19073 19904
rect 19024 19864 19030 19876
rect 19061 19873 19073 19876
rect 19107 19873 19119 19907
rect 19061 19867 19119 19873
rect 19260 19836 19288 19944
rect 19334 19932 19340 19944
rect 19392 19972 19398 19984
rect 20162 19972 20168 19984
rect 19392 19944 20168 19972
rect 19392 19932 19398 19944
rect 20162 19932 20168 19944
rect 20220 19932 20226 19984
rect 22094 19932 22100 19984
rect 22152 19972 22158 19984
rect 22152 19944 22692 19972
rect 22152 19932 22158 19944
rect 22664 19916 22692 19944
rect 23290 19932 23296 19984
rect 23348 19972 23354 19984
rect 23860 19972 23888 20003
rect 27154 20000 27160 20052
rect 27212 20040 27218 20052
rect 27341 20043 27399 20049
rect 27341 20040 27353 20043
rect 27212 20012 27353 20040
rect 27212 20000 27218 20012
rect 27341 20009 27353 20012
rect 27387 20009 27399 20043
rect 27341 20003 27399 20009
rect 23348 19944 23888 19972
rect 23348 19932 23354 19944
rect 19628 19876 19840 19904
rect 19628 19845 19656 19876
rect 18892 19808 19288 19836
rect 19613 19839 19671 19845
rect 19613 19805 19625 19839
rect 19659 19805 19671 19839
rect 19613 19799 19671 19805
rect 19702 19796 19708 19848
rect 19760 19796 19766 19848
rect 19812 19836 19840 19876
rect 19886 19864 19892 19916
rect 19944 19904 19950 19916
rect 19944 19876 20208 19904
rect 19944 19864 19950 19876
rect 19978 19836 19984 19848
rect 19812 19808 19984 19836
rect 19978 19796 19984 19808
rect 20036 19796 20042 19848
rect 20073 19839 20131 19845
rect 20073 19805 20085 19839
rect 20119 19805 20131 19839
rect 20073 19799 20131 19805
rect 18874 19728 18880 19780
rect 18932 19777 18938 19780
rect 18932 19771 18961 19777
rect 18949 19737 18961 19771
rect 18932 19731 18961 19737
rect 18932 19728 18938 19731
rect 19518 19728 19524 19780
rect 19576 19768 19582 19780
rect 20088 19768 20116 19799
rect 19576 19740 20116 19768
rect 19576 19728 19582 19740
rect 20070 19700 20076 19712
rect 18616 19672 20076 19700
rect 18417 19663 18475 19669
rect 20070 19660 20076 19672
rect 20128 19660 20134 19712
rect 20180 19700 20208 19876
rect 20346 19864 20352 19916
rect 20404 19864 20410 19916
rect 21652 19876 22508 19904
rect 20254 19796 20260 19848
rect 20312 19836 20318 19848
rect 20533 19839 20591 19845
rect 20533 19836 20545 19839
rect 20312 19808 20545 19836
rect 20312 19796 20318 19808
rect 20533 19805 20545 19808
rect 20579 19805 20591 19839
rect 20533 19799 20591 19805
rect 20548 19768 20576 19799
rect 21542 19796 21548 19848
rect 21600 19796 21606 19848
rect 21652 19845 21680 19876
rect 22480 19848 22508 19876
rect 22646 19864 22652 19916
rect 22704 19864 22710 19916
rect 22830 19864 22836 19916
rect 22888 19904 22894 19916
rect 25314 19904 25320 19916
rect 22888 19876 25320 19904
rect 22888 19864 22894 19876
rect 25314 19864 25320 19876
rect 25372 19904 25378 19916
rect 25593 19907 25651 19913
rect 25593 19904 25605 19907
rect 25372 19876 25605 19904
rect 25372 19864 25378 19876
rect 25593 19873 25605 19876
rect 25639 19904 25651 19907
rect 25958 19904 25964 19916
rect 25639 19876 25964 19904
rect 25639 19873 25651 19876
rect 25593 19867 25651 19873
rect 25958 19864 25964 19876
rect 26016 19864 26022 19916
rect 21637 19839 21695 19845
rect 21637 19805 21649 19839
rect 21683 19805 21695 19839
rect 21637 19799 21695 19805
rect 21910 19796 21916 19848
rect 21968 19796 21974 19848
rect 22002 19796 22008 19848
rect 22060 19796 22066 19848
rect 22186 19796 22192 19848
rect 22244 19836 22250 19848
rect 22281 19839 22339 19845
rect 22281 19836 22293 19839
rect 22244 19808 22293 19836
rect 22244 19796 22250 19808
rect 22281 19805 22293 19808
rect 22327 19805 22339 19839
rect 22281 19799 22339 19805
rect 22462 19796 22468 19848
rect 22520 19796 22526 19848
rect 22554 19796 22560 19848
rect 22612 19836 22618 19848
rect 22741 19839 22799 19845
rect 22741 19836 22753 19839
rect 22612 19808 22753 19836
rect 22612 19796 22618 19808
rect 22741 19805 22753 19808
rect 22787 19836 22799 19839
rect 22922 19836 22928 19848
rect 22787 19808 22928 19836
rect 22787 19805 22799 19808
rect 22741 19799 22799 19805
rect 22922 19796 22928 19808
rect 22980 19796 22986 19848
rect 23109 19839 23167 19845
rect 23109 19805 23121 19839
rect 23155 19805 23167 19839
rect 23109 19799 23167 19805
rect 21818 19768 21824 19780
rect 20548 19740 21824 19768
rect 21818 19728 21824 19740
rect 21876 19768 21882 19780
rect 21876 19740 22324 19768
rect 21876 19728 21882 19740
rect 22094 19700 22100 19712
rect 20180 19672 22100 19700
rect 22094 19660 22100 19672
rect 22152 19660 22158 19712
rect 22186 19660 22192 19712
rect 22244 19660 22250 19712
rect 22296 19700 22324 19740
rect 22370 19728 22376 19780
rect 22428 19768 22434 19780
rect 23124 19768 23152 19799
rect 23290 19796 23296 19848
rect 23348 19836 23354 19848
rect 23348 19808 23796 19836
rect 23348 19796 23354 19808
rect 22428 19740 23152 19768
rect 23569 19771 23627 19777
rect 22428 19728 22434 19740
rect 23569 19737 23581 19771
rect 23615 19768 23627 19771
rect 23658 19768 23664 19780
rect 23615 19740 23664 19768
rect 23615 19737 23627 19740
rect 23569 19731 23627 19737
rect 23658 19728 23664 19740
rect 23716 19728 23722 19780
rect 23768 19768 23796 19808
rect 23824 19771 23882 19777
rect 23824 19768 23836 19771
rect 23768 19740 23836 19768
rect 23824 19737 23836 19740
rect 23870 19737 23882 19771
rect 23824 19731 23882 19737
rect 24026 19728 24032 19780
rect 24084 19728 24090 19780
rect 25866 19728 25872 19780
rect 25924 19728 25930 19780
rect 26602 19728 26608 19780
rect 26660 19728 26666 19780
rect 24118 19700 24124 19712
rect 22296 19672 24124 19700
rect 24118 19660 24124 19672
rect 24176 19660 24182 19712
rect 1104 19610 28152 19632
rect 1104 19558 4874 19610
rect 4926 19558 4938 19610
rect 4990 19558 5002 19610
rect 5054 19558 5066 19610
rect 5118 19558 5130 19610
rect 5182 19558 28152 19610
rect 1104 19536 28152 19558
rect 1578 19456 1584 19508
rect 1636 19456 1642 19508
rect 2866 19456 2872 19508
rect 2924 19456 2930 19508
rect 3881 19499 3939 19505
rect 3881 19465 3893 19499
rect 3927 19465 3939 19499
rect 3881 19459 3939 19465
rect 5353 19499 5411 19505
rect 5353 19465 5365 19499
rect 5399 19496 5411 19499
rect 5534 19496 5540 19508
rect 5399 19468 5540 19496
rect 5399 19465 5411 19468
rect 5353 19459 5411 19465
rect 2884 19428 2912 19456
rect 3896 19428 3924 19459
rect 5534 19456 5540 19468
rect 5592 19456 5598 19508
rect 12250 19456 12256 19508
rect 12308 19496 12314 19508
rect 13630 19496 13636 19508
rect 12308 19468 13636 19496
rect 12308 19456 12314 19468
rect 13630 19456 13636 19468
rect 13688 19456 13694 19508
rect 13998 19456 14004 19508
rect 14056 19496 14062 19508
rect 15562 19496 15568 19508
rect 14056 19468 15568 19496
rect 14056 19456 14062 19468
rect 15562 19456 15568 19468
rect 15620 19456 15626 19508
rect 18506 19456 18512 19508
rect 18564 19456 18570 19508
rect 18782 19456 18788 19508
rect 18840 19496 18846 19508
rect 18840 19468 19472 19496
rect 18840 19456 18846 19468
rect 2884 19400 3096 19428
rect 3896 19400 5396 19428
rect 1394 19320 1400 19372
rect 1452 19320 1458 19372
rect 2133 19363 2191 19369
rect 2133 19329 2145 19363
rect 2179 19360 2191 19363
rect 2222 19360 2228 19372
rect 2179 19332 2228 19360
rect 2179 19329 2191 19332
rect 2133 19323 2191 19329
rect 2222 19320 2228 19332
rect 2280 19320 2286 19372
rect 2406 19320 2412 19372
rect 2464 19360 2470 19372
rect 3068 19369 3096 19400
rect 4448 19369 4476 19400
rect 2869 19363 2927 19369
rect 2869 19360 2881 19363
rect 2464 19332 2881 19360
rect 2464 19320 2470 19332
rect 2869 19329 2881 19332
rect 2915 19329 2927 19363
rect 2869 19323 2927 19329
rect 3053 19363 3111 19369
rect 3053 19329 3065 19363
rect 3099 19329 3111 19363
rect 4433 19363 4491 19369
rect 3053 19323 3111 19329
rect 3620 19332 3832 19360
rect 3620 19304 3648 19332
rect 2038 19252 2044 19304
rect 2096 19252 2102 19304
rect 2682 19252 2688 19304
rect 2740 19252 2746 19304
rect 2961 19295 3019 19301
rect 2961 19261 2973 19295
rect 3007 19292 3019 19295
rect 3421 19295 3479 19301
rect 3421 19292 3433 19295
rect 3007 19264 3433 19292
rect 3007 19261 3019 19264
rect 2961 19255 3019 19261
rect 3421 19261 3433 19264
rect 3467 19261 3479 19295
rect 3421 19255 3479 19261
rect 3513 19295 3571 19301
rect 3513 19261 3525 19295
rect 3559 19261 3571 19295
rect 3513 19255 3571 19261
rect 3528 19224 3556 19255
rect 3602 19252 3608 19304
rect 3660 19252 3666 19304
rect 3694 19252 3700 19304
rect 3752 19252 3758 19304
rect 3804 19292 3832 19332
rect 4433 19329 4445 19363
rect 4479 19329 4491 19363
rect 4433 19323 4491 19329
rect 4706 19320 4712 19372
rect 4764 19360 4770 19372
rect 5368 19369 5396 19400
rect 7852 19400 8708 19428
rect 7852 19372 7880 19400
rect 5169 19363 5227 19369
rect 5169 19360 5181 19363
rect 4764 19332 5181 19360
rect 4764 19320 4770 19332
rect 5169 19329 5181 19332
rect 5215 19329 5227 19363
rect 5169 19323 5227 19329
rect 5353 19363 5411 19369
rect 5353 19329 5365 19363
rect 5399 19329 5411 19363
rect 5353 19323 5411 19329
rect 7834 19320 7840 19372
rect 7892 19320 7898 19372
rect 8110 19320 8116 19372
rect 8168 19320 8174 19372
rect 8205 19363 8263 19369
rect 8205 19329 8217 19363
rect 8251 19360 8263 19363
rect 8386 19360 8392 19372
rect 8251 19332 8392 19360
rect 8251 19329 8263 19332
rect 8205 19323 8263 19329
rect 8386 19320 8392 19332
rect 8444 19320 8450 19372
rect 8680 19369 8708 19400
rect 14182 19388 14188 19440
rect 14240 19428 14246 19440
rect 16390 19428 16396 19440
rect 14240 19400 16396 19428
rect 14240 19388 14246 19400
rect 16390 19388 16396 19400
rect 16448 19388 16454 19440
rect 19058 19428 19064 19440
rect 18432 19400 19064 19428
rect 8665 19363 8723 19369
rect 8665 19329 8677 19363
rect 8711 19360 8723 19363
rect 8938 19360 8944 19372
rect 8711 19332 8944 19360
rect 8711 19329 8723 19332
rect 8665 19323 8723 19329
rect 8938 19320 8944 19332
rect 8996 19320 9002 19372
rect 13357 19363 13415 19369
rect 13357 19329 13369 19363
rect 13403 19329 13415 19363
rect 13357 19323 13415 19329
rect 5077 19295 5135 19301
rect 3804 19264 5028 19292
rect 4798 19224 4804 19236
rect 3528 19196 4804 19224
rect 4798 19184 4804 19196
rect 4856 19184 4862 19236
rect 5000 19224 5028 19264
rect 5077 19261 5089 19295
rect 5123 19292 5135 19295
rect 5258 19292 5264 19304
rect 5123 19264 5264 19292
rect 5123 19261 5135 19264
rect 5077 19255 5135 19261
rect 5258 19252 5264 19264
rect 5316 19252 5322 19304
rect 8573 19295 8631 19301
rect 8573 19292 8585 19295
rect 7944 19264 8585 19292
rect 7558 19224 7564 19236
rect 5000 19196 7564 19224
rect 7558 19184 7564 19196
rect 7616 19184 7622 19236
rect 7944 19168 7972 19264
rect 8573 19261 8585 19264
rect 8619 19261 8631 19295
rect 8573 19255 8631 19261
rect 13372 19236 13400 19323
rect 13722 19320 13728 19372
rect 13780 19360 13786 19372
rect 16114 19360 16120 19372
rect 13780 19332 16120 19360
rect 13780 19320 13786 19332
rect 16114 19320 16120 19332
rect 16172 19320 16178 19372
rect 18432 19369 18460 19400
rect 19058 19388 19064 19400
rect 19116 19388 19122 19440
rect 19334 19388 19340 19440
rect 19392 19388 19398 19440
rect 18417 19363 18475 19369
rect 18417 19329 18429 19363
rect 18463 19329 18475 19363
rect 18417 19323 18475 19329
rect 18690 19320 18696 19372
rect 18748 19320 18754 19372
rect 19245 19363 19303 19369
rect 19245 19329 19257 19363
rect 19291 19360 19303 19363
rect 19444 19360 19472 19468
rect 22094 19456 22100 19508
rect 22152 19496 22158 19508
rect 22554 19496 22560 19508
rect 22152 19468 22560 19496
rect 22152 19456 22158 19468
rect 22554 19456 22560 19468
rect 22612 19456 22618 19508
rect 23470 19499 23528 19505
rect 23470 19465 23482 19499
rect 23516 19496 23528 19499
rect 23566 19496 23572 19508
rect 23516 19468 23572 19496
rect 23516 19465 23528 19468
rect 23470 19459 23528 19465
rect 23566 19456 23572 19468
rect 23624 19456 23630 19508
rect 27614 19456 27620 19508
rect 27672 19456 27678 19508
rect 19702 19388 19708 19440
rect 19760 19428 19766 19440
rect 23658 19428 23664 19440
rect 19760 19400 23664 19428
rect 19760 19388 19766 19400
rect 23658 19388 23664 19400
rect 23716 19388 23722 19440
rect 19521 19363 19579 19369
rect 19521 19360 19533 19363
rect 19291 19332 19380 19360
rect 19444 19332 19533 19360
rect 19291 19329 19303 19332
rect 19245 19323 19303 19329
rect 13449 19295 13507 19301
rect 13449 19261 13461 19295
rect 13495 19261 13507 19295
rect 13449 19255 13507 19261
rect 13541 19295 13599 19301
rect 13541 19261 13553 19295
rect 13587 19261 13599 19295
rect 13541 19255 13599 19261
rect 13633 19295 13691 19301
rect 13633 19261 13645 19295
rect 13679 19292 13691 19295
rect 13814 19292 13820 19304
rect 13679 19264 13820 19292
rect 13679 19261 13691 19264
rect 13633 19255 13691 19261
rect 13354 19184 13360 19236
rect 13412 19184 13418 19236
rect 7926 19116 7932 19168
rect 7984 19116 7990 19168
rect 8202 19116 8208 19168
rect 8260 19156 8266 19168
rect 8389 19159 8447 19165
rect 8389 19156 8401 19159
rect 8260 19128 8401 19156
rect 8260 19116 8266 19128
rect 8389 19125 8401 19128
rect 8435 19125 8447 19159
rect 8389 19119 8447 19125
rect 8941 19159 8999 19165
rect 8941 19125 8953 19159
rect 8987 19156 8999 19159
rect 9674 19156 9680 19168
rect 8987 19128 9680 19156
rect 8987 19125 8999 19128
rect 8941 19119 8999 19125
rect 9674 19116 9680 19128
rect 9732 19116 9738 19168
rect 13170 19116 13176 19168
rect 13228 19116 13234 19168
rect 13262 19116 13268 19168
rect 13320 19156 13326 19168
rect 13464 19156 13492 19255
rect 13556 19224 13584 19255
rect 13814 19252 13820 19264
rect 13872 19252 13878 19304
rect 19352 19292 19380 19332
rect 19521 19329 19533 19332
rect 19567 19329 19579 19363
rect 20070 19360 20076 19372
rect 19521 19323 19579 19329
rect 19628 19332 20076 19360
rect 19628 19292 19656 19332
rect 20070 19320 20076 19332
rect 20128 19320 20134 19372
rect 22462 19320 22468 19372
rect 22520 19320 22526 19372
rect 22646 19320 22652 19372
rect 22704 19360 22710 19372
rect 22925 19363 22983 19369
rect 22925 19360 22937 19363
rect 22704 19332 22937 19360
rect 22704 19320 22710 19332
rect 22925 19329 22937 19332
rect 22971 19329 22983 19363
rect 22925 19323 22983 19329
rect 23014 19320 23020 19372
rect 23072 19360 23078 19372
rect 23290 19360 23296 19372
rect 23072 19332 23296 19360
rect 23072 19320 23078 19332
rect 23290 19320 23296 19332
rect 23348 19320 23354 19372
rect 23382 19320 23388 19372
rect 23440 19320 23446 19372
rect 23569 19363 23627 19369
rect 23569 19329 23581 19363
rect 23615 19360 23627 19363
rect 24026 19360 24032 19372
rect 23615 19332 24032 19360
rect 23615 19329 23627 19332
rect 23569 19323 23627 19329
rect 24026 19320 24032 19332
rect 24084 19320 24090 19372
rect 27798 19320 27804 19372
rect 27856 19320 27862 19372
rect 19352 19264 19656 19292
rect 15194 19224 15200 19236
rect 13556 19196 15200 19224
rect 15194 19184 15200 19196
rect 15252 19184 15258 19236
rect 19518 19184 19524 19236
rect 19576 19224 19582 19236
rect 19576 19196 22094 19224
rect 19576 19184 19582 19196
rect 13320 19128 13492 19156
rect 13320 19116 13326 19128
rect 18874 19116 18880 19168
rect 18932 19116 18938 19168
rect 19702 19116 19708 19168
rect 19760 19116 19766 19168
rect 22066 19156 22094 19196
rect 23109 19159 23167 19165
rect 23109 19156 23121 19159
rect 22066 19128 23121 19156
rect 23109 19125 23121 19128
rect 23155 19156 23167 19159
rect 23474 19156 23480 19168
rect 23155 19128 23480 19156
rect 23155 19125 23167 19128
rect 23109 19119 23167 19125
rect 23474 19116 23480 19128
rect 23532 19116 23538 19168
rect 1104 19066 28152 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 28152 19066
rect 1104 18992 28152 19014
rect 9398 18912 9404 18964
rect 9456 18952 9462 18964
rect 9493 18955 9551 18961
rect 9493 18952 9505 18955
rect 9456 18924 9505 18952
rect 9456 18912 9462 18924
rect 9493 18921 9505 18924
rect 9539 18921 9551 18955
rect 9493 18915 9551 18921
rect 13081 18955 13139 18961
rect 13081 18921 13093 18955
rect 13127 18921 13139 18955
rect 13081 18915 13139 18921
rect 2590 18844 2596 18896
rect 2648 18884 2654 18896
rect 3602 18884 3608 18896
rect 2648 18856 3608 18884
rect 2648 18844 2654 18856
rect 3602 18844 3608 18856
rect 3660 18844 3666 18896
rect 9125 18887 9183 18893
rect 9125 18853 9137 18887
rect 9171 18884 9183 18887
rect 10962 18884 10968 18896
rect 9171 18856 10968 18884
rect 9171 18853 9183 18856
rect 9125 18847 9183 18853
rect 10962 18844 10968 18856
rect 11020 18844 11026 18896
rect 13096 18884 13124 18915
rect 15102 18912 15108 18964
rect 15160 18912 15166 18964
rect 15286 18912 15292 18964
rect 15344 18912 15350 18964
rect 17773 18955 17831 18961
rect 17773 18921 17785 18955
rect 17819 18952 17831 18955
rect 19242 18952 19248 18964
rect 17819 18924 19248 18952
rect 17819 18921 17831 18924
rect 17773 18915 17831 18921
rect 15304 18884 15332 18912
rect 13096 18856 15332 18884
rect 15470 18844 15476 18896
rect 15528 18884 15534 18896
rect 17034 18884 17040 18896
rect 15528 18856 17040 18884
rect 15528 18844 15534 18856
rect 17034 18844 17040 18856
rect 17092 18844 17098 18896
rect 3620 18816 3648 18844
rect 17788 18828 17816 18915
rect 19242 18912 19248 18924
rect 19300 18912 19306 18964
rect 27798 18912 27804 18964
rect 27856 18912 27862 18964
rect 4798 18816 4804 18828
rect 3436 18788 3648 18816
rect 4540 18788 4804 18816
rect 3436 18757 3464 18788
rect 3421 18751 3479 18757
rect 3421 18717 3433 18751
rect 3467 18717 3479 18751
rect 3421 18711 3479 18717
rect 3605 18751 3663 18757
rect 3605 18717 3617 18751
rect 3651 18748 3663 18751
rect 4430 18748 4436 18760
rect 3651 18720 4436 18748
rect 3651 18717 3663 18720
rect 3605 18711 3663 18717
rect 4430 18708 4436 18720
rect 4488 18748 4494 18760
rect 4540 18757 4568 18788
rect 4798 18776 4804 18788
rect 4856 18776 4862 18828
rect 5721 18819 5779 18825
rect 5721 18785 5733 18819
rect 5767 18785 5779 18819
rect 5721 18779 5779 18785
rect 4525 18751 4583 18757
rect 4525 18748 4537 18751
rect 4488 18720 4537 18748
rect 4488 18708 4494 18720
rect 4525 18717 4537 18720
rect 4571 18717 4583 18751
rect 4525 18711 4583 18717
rect 4614 18708 4620 18760
rect 4672 18708 4678 18760
rect 5258 18708 5264 18760
rect 5316 18708 5322 18760
rect 5534 18708 5540 18760
rect 5592 18708 5598 18760
rect 5736 18748 5764 18779
rect 7926 18776 7932 18828
rect 7984 18816 7990 18828
rect 7984 18788 9168 18816
rect 7984 18776 7990 18788
rect 5905 18751 5963 18757
rect 5905 18748 5917 18751
rect 5736 18720 5917 18748
rect 5905 18717 5917 18720
rect 5951 18717 5963 18751
rect 5905 18711 5963 18717
rect 5920 18680 5948 18711
rect 6454 18708 6460 18760
rect 6512 18708 6518 18760
rect 8202 18708 8208 18760
rect 8260 18708 8266 18760
rect 8294 18708 8300 18760
rect 8352 18748 8358 18760
rect 8481 18751 8539 18757
rect 8481 18748 8493 18751
rect 8352 18720 8493 18748
rect 8352 18708 8358 18720
rect 8481 18717 8493 18720
rect 8527 18717 8539 18751
rect 8481 18711 8539 18717
rect 8938 18708 8944 18760
rect 8996 18708 9002 18760
rect 9140 18757 9168 18788
rect 13814 18776 13820 18828
rect 13872 18816 13878 18828
rect 13872 18788 14872 18816
rect 13872 18776 13878 18788
rect 9125 18751 9183 18757
rect 9125 18717 9137 18751
rect 9171 18717 9183 18751
rect 9125 18711 9183 18717
rect 9398 18708 9404 18760
rect 9456 18708 9462 18760
rect 9585 18751 9643 18757
rect 9585 18717 9597 18751
rect 9631 18717 9643 18751
rect 9585 18711 9643 18717
rect 6546 18680 6552 18692
rect 5920 18652 6552 18680
rect 6546 18640 6552 18652
rect 6604 18640 6610 18692
rect 7742 18680 7748 18692
rect 7406 18652 7748 18680
rect 7742 18640 7748 18652
rect 7800 18640 7806 18692
rect 8386 18640 8392 18692
rect 8444 18640 8450 18692
rect 9600 18680 9628 18711
rect 9674 18708 9680 18760
rect 9732 18748 9738 18760
rect 9953 18751 10011 18757
rect 9953 18748 9965 18751
rect 9732 18720 9965 18748
rect 9732 18708 9738 18720
rect 9953 18717 9965 18720
rect 9999 18717 10011 18751
rect 9953 18711 10011 18717
rect 10042 18708 10048 18760
rect 10100 18748 10106 18760
rect 10137 18751 10195 18757
rect 10137 18748 10149 18751
rect 10100 18720 10149 18748
rect 10100 18708 10106 18720
rect 10137 18717 10149 18720
rect 10183 18717 10195 18751
rect 10137 18711 10195 18717
rect 12894 18708 12900 18760
rect 12952 18708 12958 18760
rect 13078 18708 13084 18760
rect 13136 18708 13142 18760
rect 14461 18751 14519 18757
rect 14461 18717 14473 18751
rect 14507 18717 14519 18751
rect 14461 18711 14519 18717
rect 9600 18652 10088 18680
rect 3510 18572 3516 18624
rect 3568 18572 3574 18624
rect 8294 18612 8300 18624
rect 8352 18621 8358 18624
rect 8261 18584 8300 18612
rect 8294 18572 8300 18584
rect 8352 18575 8361 18621
rect 9769 18615 9827 18621
rect 9769 18581 9781 18615
rect 9815 18612 9827 18615
rect 9950 18612 9956 18624
rect 9815 18584 9956 18612
rect 9815 18581 9827 18584
rect 9769 18575 9827 18581
rect 8352 18572 8358 18575
rect 9950 18572 9956 18584
rect 10008 18572 10014 18624
rect 10060 18621 10088 18652
rect 12986 18640 12992 18692
rect 13044 18680 13050 18692
rect 14476 18680 14504 18711
rect 14642 18708 14648 18760
rect 14700 18708 14706 18760
rect 14734 18708 14740 18760
rect 14792 18708 14798 18760
rect 14844 18757 14872 18788
rect 15102 18776 15108 18828
rect 15160 18816 15166 18828
rect 17770 18816 17776 18828
rect 15160 18788 17776 18816
rect 15160 18776 15166 18788
rect 17770 18776 17776 18788
rect 17828 18776 17834 18828
rect 22741 18819 22799 18825
rect 22741 18785 22753 18819
rect 22787 18816 22799 18819
rect 22830 18816 22836 18828
rect 22787 18788 22836 18816
rect 22787 18785 22799 18788
rect 22741 18779 22799 18785
rect 22830 18776 22836 18788
rect 22888 18776 22894 18828
rect 14829 18751 14887 18757
rect 14829 18717 14841 18751
rect 14875 18717 14887 18751
rect 14829 18711 14887 18717
rect 15194 18708 15200 18760
rect 15252 18748 15258 18760
rect 15746 18748 15752 18760
rect 15252 18720 15752 18748
rect 15252 18708 15258 18720
rect 15746 18708 15752 18720
rect 15804 18708 15810 18760
rect 15838 18708 15844 18760
rect 15896 18748 15902 18760
rect 15933 18751 15991 18757
rect 15933 18748 15945 18751
rect 15896 18720 15945 18748
rect 15896 18708 15902 18720
rect 15933 18717 15945 18720
rect 15979 18748 15991 18751
rect 18506 18748 18512 18760
rect 15979 18720 18512 18748
rect 15979 18717 15991 18720
rect 15933 18711 15991 18717
rect 18506 18708 18512 18720
rect 18564 18708 18570 18760
rect 26050 18708 26056 18760
rect 26108 18708 26114 18760
rect 15212 18680 15240 18708
rect 15856 18680 15884 18708
rect 13044 18652 13400 18680
rect 14476 18652 15240 18680
rect 15304 18652 15884 18680
rect 19061 18683 19119 18689
rect 13044 18640 13050 18652
rect 13372 18624 13400 18652
rect 10045 18615 10103 18621
rect 10045 18581 10057 18615
rect 10091 18612 10103 18615
rect 10318 18612 10324 18624
rect 10091 18584 10324 18612
rect 10091 18581 10103 18584
rect 10045 18575 10103 18581
rect 10318 18572 10324 18584
rect 10376 18572 10382 18624
rect 13262 18572 13268 18624
rect 13320 18572 13326 18624
rect 13354 18572 13360 18624
rect 13412 18612 13418 18624
rect 15304 18612 15332 18652
rect 19061 18649 19073 18683
rect 19107 18680 19119 18683
rect 19334 18680 19340 18692
rect 19107 18652 19340 18680
rect 19107 18649 19119 18652
rect 19061 18643 19119 18649
rect 19334 18640 19340 18652
rect 19392 18680 19398 18692
rect 20993 18683 21051 18689
rect 20993 18680 21005 18683
rect 19392 18652 21005 18680
rect 19392 18640 19398 18652
rect 20993 18649 21005 18652
rect 21039 18649 21051 18683
rect 20993 18643 21051 18649
rect 25222 18640 25228 18692
rect 25280 18680 25286 18692
rect 26329 18683 26387 18689
rect 26329 18680 26341 18683
rect 25280 18652 26341 18680
rect 25280 18640 25286 18652
rect 26329 18649 26341 18652
rect 26375 18649 26387 18683
rect 26602 18680 26608 18692
rect 26329 18643 26387 18649
rect 26528 18652 26608 18680
rect 13412 18584 15332 18612
rect 15841 18615 15899 18621
rect 13412 18572 13418 18584
rect 15841 18581 15853 18615
rect 15887 18612 15899 18615
rect 16022 18612 16028 18624
rect 15887 18584 16028 18612
rect 15887 18581 15899 18584
rect 15841 18575 15899 18581
rect 16022 18572 16028 18584
rect 16080 18572 16086 18624
rect 24854 18572 24860 18624
rect 24912 18612 24918 18624
rect 25590 18612 25596 18624
rect 24912 18584 25596 18612
rect 24912 18572 24918 18584
rect 25590 18572 25596 18584
rect 25648 18612 25654 18624
rect 26528 18612 26556 18652
rect 26602 18640 26608 18652
rect 26660 18680 26666 18692
rect 26660 18652 26818 18680
rect 26660 18640 26666 18652
rect 25648 18584 26556 18612
rect 25648 18572 25654 18584
rect 1104 18522 28152 18544
rect 1104 18470 4874 18522
rect 4926 18470 4938 18522
rect 4990 18470 5002 18522
rect 5054 18470 5066 18522
rect 5118 18470 5130 18522
rect 5182 18470 28152 18522
rect 1104 18448 28152 18470
rect 7377 18411 7435 18417
rect 7377 18377 7389 18411
rect 7423 18408 7435 18411
rect 7926 18408 7932 18420
rect 7423 18380 7932 18408
rect 7423 18377 7435 18380
rect 7377 18371 7435 18377
rect 7926 18368 7932 18380
rect 7984 18368 7990 18420
rect 12710 18368 12716 18420
rect 12768 18408 12774 18420
rect 12989 18411 13047 18417
rect 12989 18408 13001 18411
rect 12768 18380 13001 18408
rect 12768 18368 12774 18380
rect 12989 18377 13001 18380
rect 13035 18377 13047 18411
rect 12989 18371 13047 18377
rect 13170 18368 13176 18420
rect 13228 18368 13234 18420
rect 18782 18408 18788 18420
rect 14752 18380 18788 18408
rect 4525 18343 4583 18349
rect 4525 18309 4537 18343
rect 4571 18340 4583 18343
rect 6454 18340 6460 18352
rect 4571 18312 5028 18340
rect 4571 18309 4583 18312
rect 4525 18303 4583 18309
rect 3510 18232 3516 18284
rect 3568 18232 3574 18284
rect 3694 18232 3700 18284
rect 3752 18232 3758 18284
rect 4430 18232 4436 18284
rect 4488 18232 4494 18284
rect 4614 18232 4620 18284
rect 4672 18232 4678 18284
rect 5000 18281 5028 18312
rect 6380 18312 6460 18340
rect 4985 18275 5043 18281
rect 4985 18241 4997 18275
rect 5031 18241 5043 18275
rect 4985 18235 5043 18241
rect 5258 18232 5264 18284
rect 5316 18232 5322 18284
rect 6380 18281 6408 18312
rect 6454 18300 6460 18312
rect 6512 18300 6518 18352
rect 9398 18340 9404 18352
rect 9140 18312 9404 18340
rect 6365 18275 6423 18281
rect 6365 18241 6377 18275
rect 6411 18241 6423 18275
rect 6365 18235 6423 18241
rect 6546 18232 6552 18284
rect 6604 18232 6610 18284
rect 7374 18232 7380 18284
rect 7432 18232 7438 18284
rect 7558 18232 7564 18284
rect 7616 18272 7622 18284
rect 7653 18275 7711 18281
rect 7653 18272 7665 18275
rect 7616 18244 7665 18272
rect 7616 18232 7622 18244
rect 7653 18241 7665 18244
rect 7699 18241 7711 18275
rect 7653 18235 7711 18241
rect 3970 18164 3976 18216
rect 4028 18204 4034 18216
rect 4065 18207 4123 18213
rect 4065 18204 4077 18207
rect 4028 18176 4077 18204
rect 4028 18164 4034 18176
rect 4065 18173 4077 18176
rect 4111 18173 4123 18207
rect 4065 18167 4123 18173
rect 5810 18164 5816 18216
rect 5868 18164 5874 18216
rect 6457 18207 6515 18213
rect 6457 18173 6469 18207
rect 6503 18204 6515 18207
rect 6825 18207 6883 18213
rect 6825 18204 6837 18207
rect 6503 18176 6837 18204
rect 6503 18173 6515 18176
rect 6457 18167 6515 18173
rect 6825 18173 6837 18176
rect 6871 18173 6883 18207
rect 6825 18167 6883 18173
rect 7469 18207 7527 18213
rect 7469 18173 7481 18207
rect 7515 18204 7527 18207
rect 7742 18204 7748 18216
rect 7515 18176 7748 18204
rect 7515 18173 7527 18176
rect 7469 18167 7527 18173
rect 7742 18164 7748 18176
rect 7800 18164 7806 18216
rect 7834 18164 7840 18216
rect 7892 18204 7898 18216
rect 9140 18213 9168 18312
rect 9398 18300 9404 18312
rect 9456 18300 9462 18352
rect 10965 18343 11023 18349
rect 10965 18309 10977 18343
rect 11011 18340 11023 18343
rect 14752 18340 14780 18380
rect 18782 18368 18788 18380
rect 18840 18368 18846 18420
rect 22462 18368 22468 18420
rect 22520 18408 22526 18420
rect 22738 18408 22744 18420
rect 22520 18380 22744 18408
rect 22520 18368 22526 18380
rect 22738 18368 22744 18380
rect 22796 18368 22802 18420
rect 24581 18411 24639 18417
rect 24581 18377 24593 18411
rect 24627 18408 24639 18411
rect 25130 18408 25136 18420
rect 24627 18380 25136 18408
rect 24627 18377 24639 18380
rect 24581 18371 24639 18377
rect 25130 18368 25136 18380
rect 25188 18368 25194 18420
rect 15378 18340 15384 18352
rect 11011 18312 14780 18340
rect 14844 18312 15384 18340
rect 11011 18309 11023 18312
rect 10965 18303 11023 18309
rect 9217 18275 9275 18281
rect 9217 18241 9229 18275
rect 9263 18272 9275 18275
rect 9582 18272 9588 18284
rect 9263 18244 9588 18272
rect 9263 18241 9275 18244
rect 9217 18235 9275 18241
rect 9582 18232 9588 18244
rect 9640 18232 9646 18284
rect 10042 18232 10048 18284
rect 10100 18272 10106 18284
rect 10137 18275 10195 18281
rect 10137 18272 10149 18275
rect 10100 18244 10149 18272
rect 10100 18232 10106 18244
rect 10137 18241 10149 18244
rect 10183 18241 10195 18275
rect 10137 18235 10195 18241
rect 10597 18275 10655 18281
rect 10597 18241 10609 18275
rect 10643 18272 10655 18275
rect 11054 18272 11060 18284
rect 10643 18244 11060 18272
rect 10643 18241 10655 18244
rect 10597 18235 10655 18241
rect 11054 18232 11060 18244
rect 11112 18232 11118 18284
rect 12434 18232 12440 18284
rect 12492 18272 12498 18284
rect 12805 18275 12863 18281
rect 12805 18272 12817 18275
rect 12492 18244 12817 18272
rect 12492 18232 12498 18244
rect 12805 18241 12817 18244
rect 12851 18272 12863 18275
rect 13170 18272 13176 18284
rect 12851 18244 13176 18272
rect 12851 18241 12863 18244
rect 12805 18235 12863 18241
rect 13170 18232 13176 18244
rect 13228 18232 13234 18284
rect 13262 18232 13268 18284
rect 13320 18232 13326 18284
rect 14844 18281 14872 18312
rect 15378 18300 15384 18312
rect 15436 18340 15442 18352
rect 15436 18312 16068 18340
rect 15436 18300 15442 18312
rect 13541 18275 13599 18281
rect 13541 18241 13553 18275
rect 13587 18241 13599 18275
rect 13541 18235 13599 18241
rect 14829 18275 14887 18281
rect 14829 18241 14841 18275
rect 14875 18241 14887 18275
rect 14829 18235 14887 18241
rect 9125 18207 9183 18213
rect 9125 18204 9137 18207
rect 7892 18176 9137 18204
rect 7892 18164 7898 18176
rect 9125 18173 9137 18176
rect 9171 18173 9183 18207
rect 9125 18167 9183 18173
rect 9309 18207 9367 18213
rect 9309 18173 9321 18207
rect 9355 18173 9367 18207
rect 9309 18167 9367 18173
rect 4614 18096 4620 18148
rect 4672 18136 4678 18148
rect 4672 18108 7788 18136
rect 4672 18096 4678 18108
rect 7760 18077 7788 18108
rect 8662 18096 8668 18148
rect 8720 18136 8726 18148
rect 9324 18136 9352 18167
rect 9398 18164 9404 18216
rect 9456 18164 9462 18216
rect 12066 18164 12072 18216
rect 12124 18204 12130 18216
rect 12618 18204 12624 18216
rect 12124 18176 12624 18204
rect 12124 18164 12130 18176
rect 12618 18164 12624 18176
rect 12676 18204 12682 18216
rect 12897 18207 12955 18213
rect 12897 18204 12909 18207
rect 12676 18176 12909 18204
rect 12676 18164 12682 18176
rect 12897 18173 12909 18176
rect 12943 18173 12955 18207
rect 12897 18167 12955 18173
rect 12986 18164 12992 18216
rect 13044 18204 13050 18216
rect 13449 18207 13507 18213
rect 13449 18204 13461 18207
rect 13044 18176 13461 18204
rect 13044 18164 13050 18176
rect 13449 18173 13461 18176
rect 13495 18173 13507 18207
rect 13556 18204 13584 18235
rect 15286 18232 15292 18284
rect 15344 18232 15350 18284
rect 15657 18275 15715 18281
rect 15657 18272 15669 18275
rect 15396 18244 15669 18272
rect 15304 18204 15332 18232
rect 13556 18176 15332 18204
rect 13449 18167 13507 18173
rect 9490 18136 9496 18148
rect 8720 18108 9496 18136
rect 8720 18096 8726 18108
rect 9490 18096 9496 18108
rect 9548 18096 9554 18148
rect 11882 18096 11888 18148
rect 11940 18136 11946 18148
rect 12802 18136 12808 18148
rect 11940 18108 12808 18136
rect 11940 18096 11946 18108
rect 12802 18096 12808 18108
rect 12860 18096 12866 18148
rect 13909 18139 13967 18145
rect 13909 18105 13921 18139
rect 13955 18136 13967 18139
rect 15396 18136 15424 18244
rect 15657 18241 15669 18244
rect 15703 18241 15715 18275
rect 15657 18235 15715 18241
rect 15838 18232 15844 18284
rect 15896 18232 15902 18284
rect 16040 18281 16068 18312
rect 23750 18300 23756 18352
rect 23808 18300 23814 18352
rect 16025 18275 16083 18281
rect 16025 18241 16037 18275
rect 16071 18241 16083 18275
rect 16025 18235 16083 18241
rect 16301 18275 16359 18281
rect 16301 18241 16313 18275
rect 16347 18272 16359 18275
rect 16390 18272 16396 18284
rect 16347 18244 16396 18272
rect 16347 18241 16359 18244
rect 16301 18235 16359 18241
rect 16390 18232 16396 18244
rect 16448 18232 16454 18284
rect 17770 18232 17776 18284
rect 17828 18232 17834 18284
rect 22830 18232 22836 18284
rect 22888 18232 22894 18284
rect 15470 18164 15476 18216
rect 15528 18164 15534 18216
rect 15565 18207 15623 18213
rect 15565 18173 15577 18207
rect 15611 18173 15623 18207
rect 15565 18167 15623 18173
rect 13955 18108 15424 18136
rect 15580 18136 15608 18167
rect 21910 18164 21916 18216
rect 21968 18204 21974 18216
rect 23109 18207 23167 18213
rect 23109 18204 23121 18207
rect 21968 18176 23121 18204
rect 21968 18164 21974 18176
rect 23109 18173 23121 18176
rect 23155 18173 23167 18207
rect 23109 18167 23167 18173
rect 15654 18136 15660 18148
rect 15580 18108 15660 18136
rect 13955 18105 13967 18108
rect 13909 18099 13967 18105
rect 15654 18096 15660 18108
rect 15712 18096 15718 18148
rect 16022 18096 16028 18148
rect 16080 18136 16086 18148
rect 16117 18139 16175 18145
rect 16117 18136 16129 18139
rect 16080 18108 16129 18136
rect 16080 18096 16086 18108
rect 16117 18105 16129 18108
rect 16163 18105 16175 18139
rect 16117 18099 16175 18105
rect 16209 18139 16267 18145
rect 16209 18105 16221 18139
rect 16255 18105 16267 18139
rect 16209 18099 16267 18105
rect 7745 18071 7803 18077
rect 7745 18037 7757 18071
rect 7791 18037 7803 18071
rect 7745 18031 7803 18037
rect 9585 18071 9643 18077
rect 9585 18037 9597 18071
rect 9631 18068 9643 18071
rect 9858 18068 9864 18080
rect 9631 18040 9864 18068
rect 9631 18037 9643 18040
rect 9585 18031 9643 18037
rect 9858 18028 9864 18040
rect 9916 18028 9922 18080
rect 12618 18028 12624 18080
rect 12676 18028 12682 18080
rect 14734 18028 14740 18080
rect 14792 18068 14798 18080
rect 14921 18071 14979 18077
rect 14921 18068 14933 18071
rect 14792 18040 14933 18068
rect 14792 18028 14798 18040
rect 14921 18037 14933 18040
rect 14967 18037 14979 18071
rect 14921 18031 14979 18037
rect 15010 18028 15016 18080
rect 15068 18068 15074 18080
rect 15105 18071 15163 18077
rect 15105 18068 15117 18071
rect 15068 18040 15117 18068
rect 15068 18028 15074 18040
rect 15105 18037 15117 18040
rect 15151 18068 15163 18071
rect 16224 18068 16252 18099
rect 15151 18040 16252 18068
rect 15151 18037 15163 18040
rect 15105 18031 15163 18037
rect 16482 18028 16488 18080
rect 16540 18028 16546 18080
rect 23750 18028 23756 18080
rect 23808 18068 23814 18080
rect 24854 18068 24860 18080
rect 23808 18040 24860 18068
rect 23808 18028 23814 18040
rect 24854 18028 24860 18040
rect 24912 18028 24918 18080
rect 1104 17978 28152 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 28152 17978
rect 1104 17904 28152 17926
rect 2225 17867 2283 17873
rect 2225 17833 2237 17867
rect 2271 17864 2283 17867
rect 2314 17864 2320 17876
rect 2271 17836 2320 17864
rect 2271 17833 2283 17836
rect 2225 17827 2283 17833
rect 2314 17824 2320 17836
rect 2372 17864 2378 17876
rect 2590 17864 2596 17876
rect 2372 17836 2596 17864
rect 2372 17824 2378 17836
rect 2590 17824 2596 17836
rect 2648 17824 2654 17876
rect 10965 17867 11023 17873
rect 10965 17833 10977 17867
rect 11011 17864 11023 17867
rect 11054 17864 11060 17876
rect 11011 17836 11060 17864
rect 11011 17833 11023 17836
rect 10965 17827 11023 17833
rect 11054 17824 11060 17836
rect 11112 17824 11118 17876
rect 13078 17824 13084 17876
rect 13136 17864 13142 17876
rect 13265 17867 13323 17873
rect 13265 17864 13277 17867
rect 13136 17836 13277 17864
rect 13136 17824 13142 17836
rect 13265 17833 13277 17836
rect 13311 17833 13323 17867
rect 13265 17827 13323 17833
rect 15746 17824 15752 17876
rect 15804 17864 15810 17876
rect 16761 17867 16819 17873
rect 16761 17864 16773 17867
rect 15804 17836 16773 17864
rect 15804 17824 15810 17836
rect 16761 17833 16773 17836
rect 16807 17833 16819 17867
rect 20717 17867 20775 17873
rect 20717 17864 20729 17867
rect 16761 17827 16819 17833
rect 17420 17836 20729 17864
rect 8294 17756 8300 17808
rect 8352 17796 8358 17808
rect 8941 17799 8999 17805
rect 8941 17796 8953 17799
rect 8352 17768 8953 17796
rect 8352 17756 8358 17768
rect 8941 17765 8953 17768
rect 8987 17765 8999 17799
rect 8941 17759 8999 17765
rect 9858 17756 9864 17808
rect 9916 17756 9922 17808
rect 12437 17799 12495 17805
rect 12437 17765 12449 17799
rect 12483 17796 12495 17799
rect 12483 17768 12756 17796
rect 12483 17765 12495 17768
rect 12437 17759 12495 17765
rect 9214 17688 9220 17740
rect 9272 17728 9278 17740
rect 9309 17731 9367 17737
rect 9309 17728 9321 17731
rect 9272 17700 9321 17728
rect 9272 17688 9278 17700
rect 9309 17697 9321 17700
rect 9355 17697 9367 17731
rect 9582 17728 9588 17740
rect 9309 17691 9367 17697
rect 9416 17700 9588 17728
rect 1578 17620 1584 17672
rect 1636 17660 1642 17672
rect 2317 17663 2375 17669
rect 2317 17660 2329 17663
rect 1636 17632 2329 17660
rect 1636 17620 1642 17632
rect 2317 17629 2329 17632
rect 2363 17629 2375 17663
rect 2317 17623 2375 17629
rect 7374 17620 7380 17672
rect 7432 17660 7438 17672
rect 7650 17660 7656 17672
rect 7432 17632 7656 17660
rect 7432 17620 7438 17632
rect 7650 17620 7656 17632
rect 7708 17620 7714 17672
rect 7742 17620 7748 17672
rect 7800 17620 7806 17672
rect 9122 17620 9128 17672
rect 9180 17660 9186 17672
rect 9416 17669 9444 17700
rect 9582 17688 9588 17700
rect 9640 17688 9646 17740
rect 9876 17728 9904 17756
rect 9876 17700 11284 17728
rect 9401 17663 9459 17669
rect 9401 17660 9413 17663
rect 9180 17632 9413 17660
rect 9180 17620 9186 17632
rect 9401 17629 9413 17632
rect 9447 17629 9459 17663
rect 9401 17623 9459 17629
rect 9490 17620 9496 17672
rect 9548 17660 9554 17672
rect 9861 17663 9919 17669
rect 9861 17660 9873 17663
rect 9548 17632 9873 17660
rect 9548 17620 9554 17632
rect 9861 17629 9873 17632
rect 9907 17629 9919 17663
rect 9861 17623 9919 17629
rect 10229 17663 10287 17669
rect 10229 17629 10241 17663
rect 10275 17629 10287 17663
rect 10229 17623 10287 17629
rect 8570 17552 8576 17604
rect 8628 17552 8634 17604
rect 9398 17484 9404 17536
rect 9456 17524 9462 17536
rect 10244 17524 10272 17623
rect 10318 17620 10324 17672
rect 10376 17660 10382 17672
rect 10597 17663 10655 17669
rect 10597 17660 10609 17663
rect 10376 17632 10609 17660
rect 10376 17620 10382 17632
rect 10597 17629 10609 17632
rect 10643 17629 10655 17663
rect 10597 17623 10655 17629
rect 10962 17620 10968 17672
rect 11020 17620 11026 17672
rect 11256 17669 11284 17700
rect 12158 17688 12164 17740
rect 12216 17728 12222 17740
rect 12621 17731 12679 17737
rect 12621 17728 12633 17731
rect 12216 17700 12633 17728
rect 12216 17688 12222 17700
rect 12621 17697 12633 17700
rect 12667 17697 12679 17731
rect 12728 17728 12756 17768
rect 12986 17728 12992 17740
rect 12728 17700 12992 17728
rect 12621 17691 12679 17697
rect 12986 17688 12992 17700
rect 13044 17688 13050 17740
rect 11241 17663 11299 17669
rect 11241 17629 11253 17663
rect 11287 17629 11299 17663
rect 11241 17623 11299 17629
rect 11974 17620 11980 17672
rect 12032 17660 12038 17672
rect 12250 17660 12256 17672
rect 12032 17632 12256 17660
rect 12032 17620 12038 17632
rect 12250 17620 12256 17632
rect 12308 17660 12314 17672
rect 12713 17663 12771 17669
rect 12308 17632 12572 17660
rect 12308 17620 12314 17632
rect 12544 17592 12572 17632
rect 12713 17629 12725 17663
rect 12759 17629 12771 17663
rect 13096 17660 13124 17824
rect 14829 17799 14887 17805
rect 14829 17765 14841 17799
rect 14875 17796 14887 17799
rect 15010 17796 15016 17808
rect 14875 17768 15016 17796
rect 14875 17765 14887 17768
rect 14829 17759 14887 17765
rect 15010 17756 15016 17768
rect 15068 17756 15074 17808
rect 16666 17756 16672 17808
rect 16724 17796 16730 17808
rect 17420 17796 17448 17836
rect 20717 17833 20729 17836
rect 20763 17864 20775 17867
rect 26157 17867 26215 17873
rect 26157 17864 26169 17867
rect 20763 17836 26169 17864
rect 20763 17833 20775 17836
rect 20717 17827 20775 17833
rect 19794 17796 19800 17808
rect 16724 17768 17448 17796
rect 17512 17768 19800 17796
rect 16724 17756 16730 17768
rect 12713 17623 12771 17629
rect 12912 17632 13124 17660
rect 13188 17700 13492 17728
rect 12728 17592 12756 17623
rect 12544 17564 12756 17592
rect 9456 17496 10272 17524
rect 9456 17484 9462 17496
rect 10778 17484 10784 17536
rect 10836 17524 10842 17536
rect 11149 17527 11207 17533
rect 11149 17524 11161 17527
rect 10836 17496 11161 17524
rect 10836 17484 10842 17496
rect 11149 17493 11161 17496
rect 11195 17493 11207 17527
rect 11149 17487 11207 17493
rect 11790 17484 11796 17536
rect 11848 17524 11854 17536
rect 12912 17524 12940 17632
rect 12989 17595 13047 17601
rect 12989 17561 13001 17595
rect 13035 17561 13047 17595
rect 12989 17555 13047 17561
rect 13081 17595 13139 17601
rect 13081 17561 13093 17595
rect 13127 17592 13139 17595
rect 13188 17592 13216 17700
rect 13464 17672 13492 17700
rect 14182 17688 14188 17740
rect 14240 17728 14246 17740
rect 14645 17731 14703 17737
rect 14645 17728 14657 17731
rect 14240 17700 14657 17728
rect 14240 17688 14246 17700
rect 14645 17697 14657 17700
rect 14691 17697 14703 17731
rect 16022 17728 16028 17740
rect 14645 17691 14703 17697
rect 14936 17700 16028 17728
rect 13262 17620 13268 17672
rect 13320 17660 13326 17672
rect 13357 17663 13415 17669
rect 13357 17660 13369 17663
rect 13320 17632 13369 17660
rect 13320 17620 13326 17632
rect 13357 17629 13369 17632
rect 13403 17629 13415 17663
rect 13357 17623 13415 17629
rect 13446 17620 13452 17672
rect 13504 17620 13510 17672
rect 13633 17663 13691 17669
rect 13633 17629 13645 17663
rect 13679 17660 13691 17663
rect 14826 17660 14832 17672
rect 13679 17632 14832 17660
rect 13679 17629 13691 17632
rect 13633 17623 13691 17629
rect 13648 17592 13676 17623
rect 14826 17620 14832 17632
rect 14884 17620 14890 17672
rect 14936 17669 14964 17700
rect 16022 17688 16028 17700
rect 16080 17688 16086 17740
rect 16298 17688 16304 17740
rect 16356 17728 16362 17740
rect 17512 17737 17540 17768
rect 19794 17756 19800 17768
rect 19852 17756 19858 17808
rect 20622 17756 20628 17808
rect 20680 17796 20686 17808
rect 20680 17768 22140 17796
rect 20680 17756 20686 17768
rect 17497 17731 17555 17737
rect 16356 17700 17080 17728
rect 16356 17688 16362 17700
rect 14921 17663 14979 17669
rect 14921 17629 14933 17663
rect 14967 17629 14979 17663
rect 14921 17623 14979 17629
rect 15010 17620 15016 17672
rect 15068 17620 15074 17672
rect 16390 17620 16396 17672
rect 16448 17660 16454 17672
rect 16942 17660 16948 17672
rect 16448 17632 16948 17660
rect 16448 17620 16454 17632
rect 16942 17620 16948 17632
rect 17000 17620 17006 17672
rect 17052 17669 17080 17700
rect 17497 17697 17509 17731
rect 17543 17697 17555 17731
rect 18141 17731 18199 17737
rect 18141 17728 18153 17731
rect 17497 17691 17555 17697
rect 17880 17700 18153 17728
rect 17037 17663 17095 17669
rect 17037 17629 17049 17663
rect 17083 17629 17095 17663
rect 17037 17623 17095 17629
rect 17126 17620 17132 17672
rect 17184 17620 17190 17672
rect 17770 17620 17776 17672
rect 17828 17660 17834 17672
rect 17880 17669 17908 17700
rect 18141 17697 18153 17700
rect 18187 17697 18199 17731
rect 18141 17691 18199 17697
rect 19702 17688 19708 17740
rect 19760 17728 19766 17740
rect 20349 17731 20407 17737
rect 20349 17728 20361 17731
rect 19760 17700 20361 17728
rect 19760 17688 19766 17700
rect 20349 17697 20361 17700
rect 20395 17697 20407 17731
rect 20349 17691 20407 17697
rect 20533 17731 20591 17737
rect 20533 17697 20545 17731
rect 20579 17728 20591 17731
rect 20898 17728 20904 17740
rect 20579 17700 20904 17728
rect 20579 17697 20591 17700
rect 20533 17691 20591 17697
rect 20898 17688 20904 17700
rect 20956 17688 20962 17740
rect 21177 17731 21235 17737
rect 21177 17697 21189 17731
rect 21223 17697 21235 17731
rect 22112 17728 22140 17768
rect 22186 17756 22192 17808
rect 22244 17796 22250 17808
rect 22649 17799 22707 17805
rect 22649 17796 22661 17799
rect 22244 17768 22661 17796
rect 22244 17756 22250 17768
rect 22649 17765 22661 17768
rect 22695 17765 22707 17799
rect 22649 17759 22707 17765
rect 22848 17768 24072 17796
rect 22848 17728 22876 17768
rect 22112 17700 22876 17728
rect 21177 17691 21235 17697
rect 17865 17663 17923 17669
rect 17865 17660 17877 17663
rect 17828 17632 17877 17660
rect 17828 17620 17834 17632
rect 17865 17629 17877 17632
rect 17911 17629 17923 17663
rect 17865 17623 17923 17629
rect 18049 17663 18107 17669
rect 18049 17629 18061 17663
rect 18095 17629 18107 17663
rect 18049 17623 18107 17629
rect 18325 17663 18383 17669
rect 18325 17629 18337 17663
rect 18371 17660 18383 17663
rect 18414 17660 18420 17672
rect 18371 17632 18420 17660
rect 18371 17629 18383 17632
rect 18325 17623 18383 17629
rect 15289 17595 15347 17601
rect 15289 17592 15301 17595
rect 13127 17564 13216 17592
rect 13464 17564 13676 17592
rect 14936 17564 15301 17592
rect 13127 17561 13139 17564
rect 13081 17555 13139 17561
rect 11848 17496 12940 17524
rect 13004 17524 13032 17555
rect 13464 17524 13492 17564
rect 13004 17496 13492 17524
rect 13541 17527 13599 17533
rect 11848 17484 11854 17496
rect 13541 17493 13553 17527
rect 13587 17524 13599 17527
rect 14458 17524 14464 17536
rect 13587 17496 14464 17524
rect 13587 17493 13599 17496
rect 13541 17487 13599 17493
rect 14458 17484 14464 17496
rect 14516 17484 14522 17536
rect 14550 17484 14556 17536
rect 14608 17524 14614 17536
rect 14936 17533 14964 17564
rect 15289 17561 15301 17564
rect 15335 17561 15347 17595
rect 15289 17555 15347 17561
rect 16574 17552 16580 17604
rect 16632 17592 16638 17604
rect 17144 17592 17172 17620
rect 16632 17564 17172 17592
rect 16632 17552 16638 17564
rect 17218 17552 17224 17604
rect 17276 17552 17282 17604
rect 17310 17552 17316 17604
rect 17368 17601 17374 17604
rect 17368 17595 17397 17601
rect 17385 17561 17397 17595
rect 18064 17592 18092 17623
rect 18414 17620 18420 17632
rect 18472 17620 18478 17672
rect 18601 17663 18659 17669
rect 18601 17629 18613 17663
rect 18647 17629 18659 17663
rect 18601 17623 18659 17629
rect 17368 17555 17397 17561
rect 17880 17564 18092 17592
rect 18616 17592 18644 17623
rect 18782 17620 18788 17672
rect 18840 17660 18846 17672
rect 18877 17663 18935 17669
rect 18877 17660 18889 17663
rect 18840 17632 18889 17660
rect 18840 17620 18846 17632
rect 18877 17629 18889 17632
rect 18923 17660 18935 17663
rect 19242 17660 19248 17672
rect 18923 17632 19248 17660
rect 18923 17629 18935 17632
rect 18877 17623 18935 17629
rect 19242 17620 19248 17632
rect 19300 17620 19306 17672
rect 20806 17620 20812 17672
rect 20864 17660 20870 17672
rect 21192 17660 21220 17691
rect 22572 17669 22600 17700
rect 22922 17688 22928 17740
rect 22980 17688 22986 17740
rect 23106 17688 23112 17740
rect 23164 17728 23170 17740
rect 23290 17728 23296 17740
rect 23164 17700 23296 17728
rect 23164 17688 23170 17700
rect 23290 17688 23296 17700
rect 23348 17728 23354 17740
rect 23385 17731 23443 17737
rect 23385 17728 23397 17731
rect 23348 17700 23397 17728
rect 23348 17688 23354 17700
rect 23385 17697 23397 17700
rect 23431 17697 23443 17731
rect 23385 17691 23443 17697
rect 20864 17632 21220 17660
rect 21269 17663 21327 17669
rect 20864 17620 20870 17632
rect 21269 17629 21281 17663
rect 21315 17660 21327 17663
rect 22465 17663 22523 17669
rect 22465 17660 22477 17663
rect 21315 17632 22477 17660
rect 21315 17629 21327 17632
rect 21269 17623 21327 17629
rect 22465 17629 22477 17632
rect 22511 17629 22523 17663
rect 22465 17623 22523 17629
rect 22557 17663 22615 17669
rect 22557 17629 22569 17663
rect 22603 17629 22615 17663
rect 22557 17623 22615 17629
rect 23017 17663 23075 17669
rect 23017 17629 23029 17663
rect 23063 17660 23075 17663
rect 23198 17660 23204 17672
rect 23063 17632 23204 17660
rect 23063 17629 23075 17632
rect 23017 17623 23075 17629
rect 19150 17592 19156 17604
rect 18616 17564 19156 17592
rect 17368 17552 17374 17555
rect 17880 17536 17908 17564
rect 19150 17552 19156 17564
rect 19208 17552 19214 17604
rect 20441 17595 20499 17601
rect 20441 17561 20453 17595
rect 20487 17592 20499 17595
rect 21358 17592 21364 17604
rect 20487 17564 21364 17592
rect 20487 17561 20499 17564
rect 20441 17555 20499 17561
rect 21358 17552 21364 17564
rect 21416 17552 21422 17604
rect 22480 17592 22508 17623
rect 23198 17620 23204 17632
rect 23256 17620 23262 17672
rect 23661 17663 23719 17669
rect 23661 17629 23673 17663
rect 23707 17629 23719 17663
rect 23661 17623 23719 17629
rect 23676 17592 23704 17623
rect 23842 17620 23848 17672
rect 23900 17660 23906 17672
rect 23937 17663 23995 17669
rect 23937 17660 23949 17663
rect 23900 17632 23949 17660
rect 23900 17620 23906 17632
rect 23937 17629 23949 17632
rect 23983 17629 23995 17663
rect 23937 17623 23995 17629
rect 23750 17592 23756 17604
rect 22480 17564 23756 17592
rect 23750 17552 23756 17564
rect 23808 17552 23814 17604
rect 24044 17592 24072 17768
rect 24136 17737 24164 17836
rect 26157 17833 26169 17836
rect 26203 17833 26215 17867
rect 26157 17827 26215 17833
rect 24121 17731 24179 17737
rect 24121 17697 24133 17731
rect 24167 17697 24179 17731
rect 24121 17691 24179 17697
rect 26142 17688 26148 17740
rect 26200 17728 26206 17740
rect 26421 17731 26479 17737
rect 26421 17728 26433 17731
rect 26200 17700 26433 17728
rect 26200 17688 26206 17700
rect 26421 17697 26433 17700
rect 26467 17697 26479 17731
rect 26421 17691 26479 17697
rect 24210 17620 24216 17672
rect 24268 17620 24274 17672
rect 24397 17663 24455 17669
rect 24397 17629 24409 17663
rect 24443 17660 24455 17663
rect 24486 17660 24492 17672
rect 24443 17632 24492 17660
rect 24443 17629 24455 17632
rect 24397 17623 24455 17629
rect 24486 17620 24492 17632
rect 24544 17620 24550 17672
rect 24581 17663 24639 17669
rect 24581 17629 24593 17663
rect 24627 17629 24639 17663
rect 24581 17623 24639 17629
rect 24596 17592 24624 17623
rect 24044 17564 24624 17592
rect 14921 17527 14979 17533
rect 14921 17524 14933 17527
rect 14608 17496 14933 17524
rect 14608 17484 14614 17496
rect 14921 17493 14933 17496
rect 14967 17493 14979 17527
rect 14921 17487 14979 17493
rect 16022 17484 16028 17536
rect 16080 17524 16086 17536
rect 16666 17524 16672 17536
rect 16080 17496 16672 17524
rect 16080 17484 16086 17496
rect 16666 17484 16672 17496
rect 16724 17484 16730 17536
rect 16850 17484 16856 17536
rect 16908 17484 16914 17536
rect 17862 17484 17868 17536
rect 17920 17484 17926 17536
rect 17954 17484 17960 17536
rect 18012 17484 18018 17536
rect 18509 17527 18567 17533
rect 18509 17493 18521 17527
rect 18555 17524 18567 17527
rect 18598 17524 18604 17536
rect 18555 17496 18604 17524
rect 18555 17493 18567 17496
rect 18509 17487 18567 17493
rect 18598 17484 18604 17496
rect 18656 17484 18662 17536
rect 18782 17484 18788 17536
rect 18840 17484 18846 17536
rect 20254 17484 20260 17536
rect 20312 17484 20318 17536
rect 20714 17484 20720 17536
rect 20772 17524 20778 17536
rect 20901 17527 20959 17533
rect 20901 17524 20913 17527
rect 20772 17496 20913 17524
rect 20772 17484 20778 17496
rect 20901 17493 20913 17496
rect 20947 17493 20959 17527
rect 20901 17487 20959 17493
rect 20990 17484 20996 17536
rect 21048 17524 21054 17536
rect 21542 17524 21548 17536
rect 21048 17496 21548 17524
rect 21048 17484 21054 17496
rect 21542 17484 21548 17496
rect 21600 17524 21606 17536
rect 23198 17524 23204 17536
rect 21600 17496 23204 17524
rect 21600 17484 21606 17496
rect 23198 17484 23204 17496
rect 23256 17484 23262 17536
rect 24394 17484 24400 17536
rect 24452 17524 24458 17536
rect 24489 17527 24547 17533
rect 24489 17524 24501 17527
rect 24452 17496 24501 17524
rect 24452 17484 24458 17496
rect 24489 17493 24501 17496
rect 24535 17493 24547 17527
rect 24596 17524 24624 17564
rect 24854 17552 24860 17604
rect 24912 17592 24918 17604
rect 24912 17564 24978 17592
rect 24912 17552 24918 17564
rect 24673 17527 24731 17533
rect 24673 17524 24685 17527
rect 24596 17496 24685 17524
rect 24489 17487 24547 17493
rect 24673 17493 24685 17496
rect 24719 17524 24731 17527
rect 24762 17524 24768 17536
rect 24719 17496 24768 17524
rect 24719 17493 24731 17496
rect 24673 17487 24731 17493
rect 24762 17484 24768 17496
rect 24820 17484 24826 17536
rect 1104 17434 28152 17456
rect 1104 17382 4874 17434
rect 4926 17382 4938 17434
rect 4990 17382 5002 17434
rect 5054 17382 5066 17434
rect 5118 17382 5130 17434
rect 5182 17382 28152 17434
rect 1104 17360 28152 17382
rect 2682 17320 2688 17332
rect 2608 17292 2688 17320
rect 1857 17255 1915 17261
rect 1857 17221 1869 17255
rect 1903 17252 1915 17255
rect 2038 17252 2044 17264
rect 1903 17224 2044 17252
rect 1903 17221 1915 17224
rect 1857 17215 1915 17221
rect 2038 17212 2044 17224
rect 2096 17252 2102 17264
rect 2498 17252 2504 17264
rect 2096 17224 2504 17252
rect 2096 17212 2102 17224
rect 2498 17212 2504 17224
rect 2556 17212 2562 17264
rect 842 17144 848 17196
rect 900 17184 906 17196
rect 1489 17187 1547 17193
rect 1489 17184 1501 17187
rect 900 17156 1501 17184
rect 900 17144 906 17156
rect 1489 17153 1501 17156
rect 1535 17153 1547 17187
rect 2608 17170 2636 17292
rect 2682 17280 2688 17292
rect 2740 17320 2746 17332
rect 15010 17320 15016 17332
rect 2740 17292 3372 17320
rect 2740 17280 2746 17292
rect 3053 17255 3111 17261
rect 3053 17221 3065 17255
rect 3099 17252 3111 17255
rect 3234 17252 3240 17264
rect 3099 17224 3240 17252
rect 3099 17221 3111 17224
rect 3053 17215 3111 17221
rect 3234 17212 3240 17224
rect 3292 17212 3298 17264
rect 3344 17193 3372 17292
rect 12084 17292 15016 17320
rect 10594 17212 10600 17264
rect 10652 17252 10658 17264
rect 12084 17252 12112 17292
rect 15010 17280 15016 17292
rect 15068 17280 15074 17332
rect 16393 17323 16451 17329
rect 16393 17289 16405 17323
rect 16439 17320 16451 17323
rect 16574 17320 16580 17332
rect 16439 17292 16580 17320
rect 16439 17289 16451 17292
rect 16393 17283 16451 17289
rect 16574 17280 16580 17292
rect 16632 17280 16638 17332
rect 16761 17323 16819 17329
rect 16761 17289 16773 17323
rect 16807 17320 16819 17323
rect 17310 17320 17316 17332
rect 16807 17292 17316 17320
rect 16807 17289 16819 17292
rect 16761 17283 16819 17289
rect 17310 17280 17316 17292
rect 17368 17280 17374 17332
rect 18598 17280 18604 17332
rect 18656 17320 18662 17332
rect 19889 17323 19947 17329
rect 19889 17320 19901 17323
rect 18656 17292 19901 17320
rect 18656 17280 18662 17292
rect 19889 17289 19901 17292
rect 19935 17289 19947 17323
rect 19889 17283 19947 17289
rect 20530 17280 20536 17332
rect 20588 17280 20594 17332
rect 21910 17280 21916 17332
rect 21968 17280 21974 17332
rect 23937 17323 23995 17329
rect 23937 17289 23949 17323
rect 23983 17320 23995 17323
rect 24210 17320 24216 17332
rect 23983 17292 24216 17320
rect 23983 17289 23995 17292
rect 23937 17283 23995 17289
rect 24210 17280 24216 17292
rect 24268 17280 24274 17332
rect 12802 17252 12808 17264
rect 10652 17224 12112 17252
rect 10652 17212 10658 17224
rect 3145 17187 3203 17193
rect 1489 17147 1547 17153
rect 3145 17153 3157 17187
rect 3191 17153 3203 17187
rect 3145 17147 3203 17153
rect 3329 17187 3387 17193
rect 3329 17153 3341 17187
rect 3375 17153 3387 17187
rect 3329 17147 3387 17153
rect 2225 17119 2283 17125
rect 2225 17085 2237 17119
rect 2271 17085 2283 17119
rect 2225 17079 2283 17085
rect 2240 17048 2268 17079
rect 2406 17048 2412 17060
rect 2240 17020 2412 17048
rect 2406 17008 2412 17020
rect 2464 17048 2470 17060
rect 3160 17048 3188 17147
rect 3786 17144 3792 17196
rect 3844 17144 3850 17196
rect 3970 17144 3976 17196
rect 4028 17144 4034 17196
rect 7282 17144 7288 17196
rect 7340 17144 7346 17196
rect 8018 17144 8024 17196
rect 8076 17144 8082 17196
rect 8570 17144 8576 17196
rect 8628 17144 8634 17196
rect 9858 17144 9864 17196
rect 9916 17144 9922 17196
rect 9950 17144 9956 17196
rect 10008 17184 10014 17196
rect 10045 17187 10103 17193
rect 10045 17184 10057 17187
rect 10008 17156 10057 17184
rect 10008 17144 10014 17156
rect 10045 17153 10057 17156
rect 10091 17184 10103 17187
rect 10778 17184 10784 17196
rect 10091 17156 10784 17184
rect 10091 17153 10103 17156
rect 10045 17147 10103 17153
rect 10778 17144 10784 17156
rect 10836 17144 10842 17196
rect 11790 17144 11796 17196
rect 11848 17144 11854 17196
rect 11882 17144 11888 17196
rect 11940 17144 11946 17196
rect 11974 17144 11980 17196
rect 12032 17144 12038 17196
rect 5626 17076 5632 17128
rect 5684 17116 5690 17128
rect 6365 17119 6423 17125
rect 6365 17116 6377 17119
rect 5684 17088 6377 17116
rect 5684 17076 5690 17088
rect 6365 17085 6377 17088
rect 6411 17085 6423 17119
rect 6365 17079 6423 17085
rect 6914 17076 6920 17128
rect 6972 17116 6978 17128
rect 7377 17119 7435 17125
rect 7377 17116 7389 17119
rect 6972 17088 7389 17116
rect 6972 17076 6978 17088
rect 7377 17085 7389 17088
rect 7423 17085 7435 17119
rect 7377 17079 7435 17085
rect 10870 17076 10876 17128
rect 10928 17076 10934 17128
rect 12084 17116 12112 17224
rect 12268 17224 12808 17252
rect 12161 17187 12219 17193
rect 12161 17153 12173 17187
rect 12207 17184 12219 17187
rect 12268 17184 12296 17224
rect 12802 17212 12808 17224
rect 12860 17212 12866 17264
rect 14458 17212 14464 17264
rect 14516 17252 14522 17264
rect 14516 17224 14872 17252
rect 14516 17212 14522 17224
rect 12207 17156 12296 17184
rect 12207 17153 12219 17156
rect 12161 17147 12219 17153
rect 13630 17144 13636 17196
rect 13688 17144 13694 17196
rect 14550 17144 14556 17196
rect 14608 17144 14614 17196
rect 14734 17144 14740 17196
rect 14792 17144 14798 17196
rect 14844 17184 14872 17224
rect 17954 17212 17960 17264
rect 18012 17212 18018 17264
rect 20073 17255 20131 17261
rect 20073 17252 20085 17255
rect 19260 17224 20085 17252
rect 15749 17187 15807 17193
rect 15749 17184 15761 17187
rect 14844 17156 15761 17184
rect 15749 17153 15761 17156
rect 15795 17153 15807 17187
rect 15749 17147 15807 17153
rect 15838 17144 15844 17196
rect 15896 17184 15902 17196
rect 15933 17187 15991 17193
rect 15933 17184 15945 17187
rect 15896 17156 15945 17184
rect 15896 17144 15902 17156
rect 15933 17153 15945 17156
rect 15979 17153 15991 17187
rect 15933 17147 15991 17153
rect 16022 17144 16028 17196
rect 16080 17182 16086 17196
rect 16117 17187 16175 17193
rect 16117 17182 16129 17187
rect 16080 17154 16129 17182
rect 16080 17144 16086 17154
rect 16117 17153 16129 17154
rect 16163 17153 16175 17187
rect 16117 17147 16175 17153
rect 16206 17144 16212 17196
rect 16264 17144 16270 17196
rect 16298 17144 16304 17196
rect 16356 17184 16362 17196
rect 16485 17187 16543 17193
rect 16356 17182 16436 17184
rect 16485 17182 16497 17187
rect 16356 17156 16497 17182
rect 16356 17144 16362 17156
rect 16408 17154 16497 17156
rect 16485 17153 16497 17154
rect 16531 17153 16543 17187
rect 16485 17147 16543 17153
rect 16666 17144 16672 17196
rect 16724 17144 16730 17196
rect 16942 17144 16948 17196
rect 17000 17144 17006 17196
rect 17126 17144 17132 17196
rect 17184 17184 17190 17196
rect 17221 17187 17279 17193
rect 17221 17184 17233 17187
rect 17184 17156 17233 17184
rect 17184 17144 17190 17156
rect 17221 17153 17233 17156
rect 17267 17153 17279 17187
rect 17221 17147 17279 17153
rect 17678 17144 17684 17196
rect 17736 17144 17742 17196
rect 19058 17144 19064 17196
rect 19116 17144 19122 17196
rect 19260 17184 19288 17224
rect 20073 17221 20085 17224
rect 20119 17221 20131 17255
rect 24029 17255 24087 17261
rect 24029 17252 24041 17255
rect 20073 17215 20131 17221
rect 20180 17224 20944 17252
rect 19168 17156 19288 17184
rect 19705 17187 19763 17193
rect 12253 17119 12311 17125
rect 12253 17116 12265 17119
rect 12084 17088 12265 17116
rect 12253 17085 12265 17088
rect 12299 17085 12311 17119
rect 12253 17079 12311 17085
rect 12529 17119 12587 17125
rect 12529 17085 12541 17119
rect 12575 17116 12587 17119
rect 13538 17116 13544 17128
rect 12575 17088 13544 17116
rect 12575 17085 12587 17088
rect 12529 17079 12587 17085
rect 13538 17076 13544 17088
rect 13596 17076 13602 17128
rect 13906 17076 13912 17128
rect 13964 17116 13970 17128
rect 15013 17119 15071 17125
rect 15013 17116 15025 17119
rect 13964 17088 15025 17116
rect 13964 17076 13970 17088
rect 15013 17085 15025 17088
rect 15059 17085 15071 17119
rect 15013 17079 15071 17085
rect 15289 17119 15347 17125
rect 15289 17085 15301 17119
rect 15335 17116 15347 17119
rect 15335 17088 16620 17116
rect 15335 17085 15347 17088
rect 15289 17079 15347 17085
rect 2464 17020 3188 17048
rect 6825 17051 6883 17057
rect 2464 17008 2470 17020
rect 6825 17017 6837 17051
rect 6871 17048 6883 17051
rect 8018 17048 8024 17060
rect 6871 17020 8024 17048
rect 6871 17017 6883 17020
rect 6825 17011 6883 17017
rect 8018 17008 8024 17020
rect 8076 17008 8082 17060
rect 11701 17051 11759 17057
rect 11701 17017 11713 17051
rect 11747 17048 11759 17051
rect 14921 17051 14979 17057
rect 11747 17020 12112 17048
rect 11747 17017 11759 17020
rect 11701 17011 11759 17017
rect 2958 16940 2964 16992
rect 3016 16980 3022 16992
rect 3329 16983 3387 16989
rect 3329 16980 3341 16983
rect 3016 16952 3341 16980
rect 3016 16940 3022 16952
rect 3329 16949 3341 16952
rect 3375 16949 3387 16983
rect 3329 16943 3387 16949
rect 3878 16940 3884 16992
rect 3936 16940 3942 16992
rect 9493 16983 9551 16989
rect 9493 16949 9505 16983
rect 9539 16980 9551 16983
rect 9766 16980 9772 16992
rect 9539 16952 9772 16980
rect 9539 16949 9551 16952
rect 9493 16943 9551 16949
rect 9766 16940 9772 16952
rect 9824 16940 9830 16992
rect 12084 16980 12112 17020
rect 14921 17017 14933 17051
rect 14967 17048 14979 17051
rect 16209 17051 16267 17057
rect 16209 17048 16221 17051
rect 14967 17020 16221 17048
rect 14967 17017 14979 17020
rect 14921 17011 14979 17017
rect 16209 17017 16221 17020
rect 16255 17017 16267 17051
rect 16209 17011 16267 17017
rect 12894 16980 12900 16992
rect 12084 16952 12900 16980
rect 12894 16940 12900 16952
rect 12952 16940 12958 16992
rect 13262 16940 13268 16992
rect 13320 16980 13326 16992
rect 13814 16980 13820 16992
rect 13320 16952 13820 16980
rect 13320 16940 13326 16952
rect 13814 16940 13820 16952
rect 13872 16980 13878 16992
rect 14001 16983 14059 16989
rect 14001 16980 14013 16983
rect 13872 16952 14013 16980
rect 13872 16940 13878 16952
rect 14001 16949 14013 16952
rect 14047 16949 14059 16983
rect 14001 16943 14059 16949
rect 14826 16940 14832 16992
rect 14884 16940 14890 16992
rect 15378 16940 15384 16992
rect 15436 16940 15442 16992
rect 15654 16940 15660 16992
rect 15712 16940 15718 16992
rect 15841 16983 15899 16989
rect 15841 16949 15853 16983
rect 15887 16980 15899 16983
rect 16482 16980 16488 16992
rect 15887 16952 16488 16980
rect 15887 16949 15899 16952
rect 15841 16943 15899 16949
rect 16482 16940 16488 16952
rect 16540 16940 16546 16992
rect 16592 16980 16620 17088
rect 17034 17076 17040 17128
rect 17092 17076 17098 17128
rect 17310 17076 17316 17128
rect 17368 17116 17374 17128
rect 19168 17116 19196 17156
rect 19705 17153 19717 17187
rect 19751 17184 19763 17187
rect 19981 17187 20039 17193
rect 19981 17184 19993 17187
rect 19751 17156 19993 17184
rect 19751 17153 19763 17156
rect 19705 17147 19763 17153
rect 19981 17153 19993 17156
rect 20027 17184 20039 17187
rect 20180 17184 20208 17224
rect 20916 17196 20944 17224
rect 23400 17224 24041 17252
rect 20027 17156 20208 17184
rect 20027 17153 20039 17156
rect 19981 17147 20039 17153
rect 20254 17144 20260 17196
rect 20312 17144 20318 17196
rect 20346 17144 20352 17196
rect 20404 17144 20410 17196
rect 20622 17144 20628 17196
rect 20680 17144 20686 17196
rect 20806 17144 20812 17196
rect 20864 17144 20870 17196
rect 20898 17144 20904 17196
rect 20956 17144 20962 17196
rect 20993 17187 21051 17193
rect 20993 17153 21005 17187
rect 21039 17153 21051 17187
rect 20993 17147 21051 17153
rect 21100 17156 21496 17184
rect 17368 17088 19196 17116
rect 17368 17076 17374 17088
rect 20530 17076 20536 17128
rect 20588 17116 20594 17128
rect 21008 17116 21036 17147
rect 20588 17088 21036 17116
rect 20588 17076 20594 17088
rect 21100 17048 21128 17156
rect 21269 17119 21327 17125
rect 21269 17085 21281 17119
rect 21315 17085 21327 17119
rect 21468 17116 21496 17156
rect 21542 17144 21548 17196
rect 21600 17144 21606 17196
rect 21818 17144 21824 17196
rect 21876 17144 21882 17196
rect 22005 17187 22063 17193
rect 22005 17153 22017 17187
rect 22051 17153 22063 17187
rect 22005 17147 22063 17153
rect 22020 17116 22048 17147
rect 22094 17144 22100 17196
rect 22152 17184 22158 17196
rect 23198 17184 23204 17196
rect 22152 17156 23204 17184
rect 22152 17144 22158 17156
rect 23198 17144 23204 17156
rect 23256 17144 23262 17196
rect 23400 17193 23428 17224
rect 24029 17221 24041 17224
rect 24075 17221 24087 17255
rect 24029 17215 24087 17221
rect 24394 17212 24400 17264
rect 24452 17212 24458 17264
rect 23385 17187 23443 17193
rect 23385 17153 23397 17187
rect 23431 17153 23443 17187
rect 23385 17147 23443 17153
rect 23474 17144 23480 17196
rect 23532 17144 23538 17196
rect 23750 17144 23756 17196
rect 23808 17144 23814 17196
rect 24213 17187 24271 17193
rect 24213 17153 24225 17187
rect 24259 17153 24271 17187
rect 24213 17147 24271 17153
rect 21468 17088 22048 17116
rect 23569 17119 23627 17125
rect 21269 17079 21327 17085
rect 23569 17085 23581 17119
rect 23615 17116 23627 17119
rect 23658 17116 23664 17128
rect 23615 17088 23664 17116
rect 23615 17085 23627 17088
rect 23569 17079 23627 17085
rect 19812 17020 21128 17048
rect 21177 17051 21235 17057
rect 16945 16983 17003 16989
rect 16945 16980 16957 16983
rect 16592 16952 16957 16980
rect 16945 16949 16957 16952
rect 16991 16949 17003 16983
rect 16945 16943 17003 16949
rect 17405 16983 17463 16989
rect 17405 16949 17417 16983
rect 17451 16980 17463 16983
rect 19812 16980 19840 17020
rect 21177 17017 21189 17051
rect 21223 17048 21235 17051
rect 21284 17048 21312 17079
rect 23658 17076 23664 17088
rect 23716 17116 23722 17128
rect 23934 17116 23940 17128
rect 23716 17088 23940 17116
rect 23716 17076 23722 17088
rect 23934 17076 23940 17088
rect 23992 17076 23998 17128
rect 24228 17116 24256 17147
rect 24486 17144 24492 17196
rect 24544 17184 24550 17196
rect 24673 17187 24731 17193
rect 24673 17184 24685 17187
rect 24544 17156 24685 17184
rect 24544 17144 24550 17156
rect 24673 17153 24685 17156
rect 24719 17153 24731 17187
rect 24673 17147 24731 17153
rect 24762 17144 24768 17196
rect 24820 17144 24826 17196
rect 24228 17088 24532 17116
rect 21223 17020 21312 17048
rect 21223 17017 21235 17020
rect 21177 17011 21235 17017
rect 22922 17008 22928 17060
rect 22980 17048 22986 17060
rect 24228 17048 24256 17088
rect 24504 17057 24532 17088
rect 22980 17020 24256 17048
rect 24489 17051 24547 17057
rect 22980 17008 22986 17020
rect 24489 17017 24501 17051
rect 24535 17017 24547 17051
rect 24489 17011 24547 17017
rect 17451 16952 19840 16980
rect 17451 16949 17463 16952
rect 17405 16943 17463 16949
rect 19886 16940 19892 16992
rect 19944 16980 19950 16992
rect 20073 16983 20131 16989
rect 20073 16980 20085 16983
rect 19944 16952 20085 16980
rect 19944 16940 19950 16952
rect 20073 16949 20085 16952
rect 20119 16949 20131 16983
rect 20073 16943 20131 16949
rect 20806 16940 20812 16992
rect 20864 16980 20870 16992
rect 21361 16983 21419 16989
rect 21361 16980 21373 16983
rect 20864 16952 21373 16980
rect 20864 16940 20870 16952
rect 21361 16949 21373 16952
rect 21407 16949 21419 16983
rect 21361 16943 21419 16949
rect 21450 16940 21456 16992
rect 21508 16940 21514 16992
rect 1104 16890 28152 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 28152 16890
rect 1104 16816 28152 16838
rect 2406 16736 2412 16788
rect 2464 16736 2470 16788
rect 7745 16779 7803 16785
rect 7745 16745 7757 16779
rect 7791 16776 7803 16779
rect 7834 16776 7840 16788
rect 7791 16748 7840 16776
rect 7791 16745 7803 16748
rect 7745 16739 7803 16745
rect 7834 16736 7840 16748
rect 7892 16736 7898 16788
rect 9309 16779 9367 16785
rect 9309 16745 9321 16779
rect 9355 16776 9367 16779
rect 9398 16776 9404 16788
rect 9355 16748 9404 16776
rect 9355 16745 9367 16748
rect 9309 16739 9367 16745
rect 9398 16736 9404 16748
rect 9456 16736 9462 16788
rect 13446 16736 13452 16788
rect 13504 16736 13510 16788
rect 13630 16736 13636 16788
rect 13688 16776 13694 16788
rect 17405 16779 17463 16785
rect 13688 16748 15976 16776
rect 13688 16736 13694 16748
rect 4614 16708 4620 16720
rect 1964 16680 3188 16708
rect 1964 16649 1992 16680
rect 3160 16652 3188 16680
rect 3344 16680 4620 16708
rect 1949 16643 2007 16649
rect 1949 16609 1961 16643
rect 1995 16609 2007 16643
rect 2225 16643 2283 16649
rect 2225 16640 2237 16643
rect 1949 16603 2007 16609
rect 2148 16612 2237 16640
rect 1857 16575 1915 16581
rect 1857 16541 1869 16575
rect 1903 16572 1915 16575
rect 2038 16572 2044 16584
rect 1903 16544 2044 16572
rect 1903 16541 1915 16544
rect 1857 16535 1915 16541
rect 2038 16532 2044 16544
rect 2096 16532 2102 16584
rect 2148 16572 2176 16612
rect 2225 16609 2237 16612
rect 2271 16640 2283 16643
rect 2314 16640 2320 16652
rect 2271 16612 2320 16640
rect 2271 16609 2283 16612
rect 2225 16603 2283 16609
rect 2314 16600 2320 16612
rect 2372 16600 2378 16652
rect 3142 16600 3148 16652
rect 3200 16600 3206 16652
rect 3234 16600 3240 16652
rect 3292 16600 3298 16652
rect 2148 16571 2360 16572
rect 2148 16565 2375 16571
rect 2148 16544 2329 16565
rect 2317 16531 2329 16544
rect 2363 16531 2375 16565
rect 2498 16532 2504 16584
rect 2556 16532 2562 16584
rect 2958 16532 2964 16584
rect 3016 16532 3022 16584
rect 3053 16575 3111 16581
rect 3053 16541 3065 16575
rect 3099 16572 3111 16575
rect 3344 16572 3372 16680
rect 4614 16668 4620 16680
rect 4672 16708 4678 16720
rect 5350 16708 5356 16720
rect 4672 16680 5356 16708
rect 4672 16668 4678 16680
rect 5350 16668 5356 16680
rect 5408 16668 5414 16720
rect 10870 16668 10876 16720
rect 10928 16708 10934 16720
rect 15838 16708 15844 16720
rect 10928 16680 15844 16708
rect 10928 16668 10934 16680
rect 15838 16668 15844 16680
rect 15896 16668 15902 16720
rect 15948 16708 15976 16748
rect 17405 16745 17417 16779
rect 17451 16776 17463 16779
rect 17494 16776 17500 16788
rect 17451 16748 17500 16776
rect 17451 16745 17463 16748
rect 17405 16739 17463 16745
rect 17494 16736 17500 16748
rect 17552 16736 17558 16788
rect 17727 16779 17785 16785
rect 17727 16776 17739 16779
rect 17604 16748 17739 16776
rect 16390 16708 16396 16720
rect 15948 16680 16396 16708
rect 16390 16668 16396 16680
rect 16448 16668 16454 16720
rect 17310 16708 17316 16720
rect 17144 16680 17316 16708
rect 3421 16643 3479 16649
rect 3421 16609 3433 16643
rect 3467 16640 3479 16643
rect 3786 16640 3792 16652
rect 3467 16612 3792 16640
rect 3467 16609 3479 16612
rect 3421 16603 3479 16609
rect 3786 16600 3792 16612
rect 3844 16640 3850 16652
rect 4065 16643 4123 16649
rect 4065 16640 4077 16643
rect 3844 16612 4077 16640
rect 3844 16600 3850 16612
rect 4065 16609 4077 16612
rect 4111 16609 4123 16643
rect 9766 16640 9772 16652
rect 4065 16603 4123 16609
rect 5092 16612 5488 16640
rect 3099 16544 3372 16572
rect 3099 16541 3111 16544
rect 3053 16535 3111 16541
rect 3970 16532 3976 16584
rect 4028 16572 4034 16584
rect 4157 16575 4215 16581
rect 4157 16572 4169 16575
rect 4028 16544 4169 16572
rect 4028 16532 4034 16544
rect 4157 16541 4169 16544
rect 4203 16541 4215 16575
rect 4157 16535 4215 16541
rect 4522 16532 4528 16584
rect 4580 16572 4586 16584
rect 5092 16581 5120 16612
rect 5460 16581 5488 16612
rect 9324 16612 9772 16640
rect 5077 16575 5135 16581
rect 5077 16572 5089 16575
rect 4580 16544 5089 16572
rect 4580 16532 4586 16544
rect 5077 16541 5089 16544
rect 5123 16541 5135 16575
rect 5077 16535 5135 16541
rect 5261 16575 5319 16581
rect 5261 16541 5273 16575
rect 5307 16541 5319 16575
rect 5261 16535 5319 16541
rect 5445 16575 5503 16581
rect 5445 16541 5457 16575
rect 5491 16541 5503 16575
rect 5445 16535 5503 16541
rect 2317 16525 2375 16531
rect 5276 16504 5304 16535
rect 5810 16532 5816 16584
rect 5868 16572 5874 16584
rect 5997 16575 6055 16581
rect 5997 16572 6009 16575
rect 5868 16544 6009 16572
rect 5868 16532 5874 16544
rect 5997 16541 6009 16544
rect 6043 16541 6055 16575
rect 5997 16535 6055 16541
rect 8018 16532 8024 16584
rect 8076 16532 8082 16584
rect 8478 16532 8484 16584
rect 8536 16572 8542 16584
rect 8573 16575 8631 16581
rect 8573 16572 8585 16575
rect 8536 16544 8585 16572
rect 8536 16532 8542 16544
rect 8573 16541 8585 16544
rect 8619 16541 8631 16575
rect 8573 16535 8631 16541
rect 9030 16532 9036 16584
rect 9088 16572 9094 16584
rect 9324 16581 9352 16612
rect 9766 16600 9772 16612
rect 9824 16600 9830 16652
rect 12618 16600 12624 16652
rect 12676 16640 12682 16652
rect 12989 16643 13047 16649
rect 12989 16640 13001 16643
rect 12676 16612 13001 16640
rect 12676 16600 12682 16612
rect 12989 16609 13001 16612
rect 13035 16609 13047 16643
rect 12989 16603 13047 16609
rect 13081 16643 13139 16649
rect 13081 16609 13093 16643
rect 13127 16640 13139 16643
rect 13354 16640 13360 16652
rect 13127 16612 13360 16640
rect 13127 16609 13139 16612
rect 13081 16603 13139 16609
rect 13354 16600 13360 16612
rect 13412 16600 13418 16652
rect 15378 16600 15384 16652
rect 15436 16640 15442 16652
rect 17144 16640 17172 16680
rect 17310 16668 17316 16680
rect 17368 16668 17374 16720
rect 15436 16612 17172 16640
rect 17221 16643 17279 16649
rect 15436 16600 15442 16612
rect 17221 16609 17233 16643
rect 17267 16640 17279 16643
rect 17604 16640 17632 16748
rect 17727 16745 17739 16748
rect 17773 16776 17785 16779
rect 17862 16776 17868 16788
rect 17773 16748 17868 16776
rect 17773 16745 17785 16748
rect 17727 16739 17785 16745
rect 17862 16736 17868 16748
rect 17920 16776 17926 16788
rect 18141 16779 18199 16785
rect 18141 16776 18153 16779
rect 17920 16748 18153 16776
rect 17920 16736 17926 16748
rect 18141 16745 18153 16748
rect 18187 16745 18199 16779
rect 18782 16776 18788 16788
rect 18141 16739 18199 16745
rect 18248 16748 18788 16776
rect 18248 16708 18276 16748
rect 18782 16736 18788 16748
rect 18840 16736 18846 16788
rect 19794 16736 19800 16788
rect 19852 16776 19858 16788
rect 22094 16776 22100 16788
rect 19852 16748 22100 16776
rect 19852 16736 19858 16748
rect 22094 16736 22100 16748
rect 22152 16736 22158 16788
rect 25498 16736 25504 16788
rect 25556 16776 25562 16788
rect 26329 16779 26387 16785
rect 26329 16776 26341 16779
rect 25556 16748 26341 16776
rect 25556 16736 25562 16748
rect 26329 16745 26341 16748
rect 26375 16745 26387 16779
rect 26329 16739 26387 16745
rect 17267 16612 17448 16640
rect 17267 16609 17279 16612
rect 17221 16603 17279 16609
rect 9125 16575 9183 16581
rect 9125 16572 9137 16575
rect 9088 16544 9137 16572
rect 9088 16532 9094 16544
rect 9125 16541 9137 16544
rect 9171 16541 9183 16575
rect 9125 16535 9183 16541
rect 9309 16575 9367 16581
rect 9309 16541 9321 16575
rect 9355 16541 9367 16575
rect 9309 16535 9367 16541
rect 12069 16575 12127 16581
rect 12069 16541 12081 16575
rect 12115 16572 12127 16575
rect 12158 16572 12164 16584
rect 12115 16544 12164 16572
rect 12115 16541 12127 16544
rect 12069 16535 12127 16541
rect 12158 16532 12164 16544
rect 12216 16532 12222 16584
rect 12250 16532 12256 16584
rect 12308 16532 12314 16584
rect 12437 16575 12495 16581
rect 12437 16541 12449 16575
rect 12483 16541 12495 16575
rect 12437 16535 12495 16541
rect 12713 16575 12771 16581
rect 12713 16541 12725 16575
rect 12759 16541 12771 16575
rect 12713 16535 12771 16541
rect 5828 16504 5856 16532
rect 5276 16476 5856 16504
rect 6920 16516 6972 16522
rect 7558 16464 7564 16516
rect 7616 16504 7622 16516
rect 7745 16507 7803 16513
rect 7745 16504 7757 16507
rect 7616 16476 7757 16504
rect 7616 16464 7622 16476
rect 7745 16473 7757 16476
rect 7791 16473 7803 16507
rect 7745 16467 7803 16473
rect 8294 16464 8300 16516
rect 8352 16504 8358 16516
rect 8389 16507 8447 16513
rect 8389 16504 8401 16507
rect 8352 16476 8401 16504
rect 8352 16464 8358 16476
rect 8389 16473 8401 16476
rect 8435 16473 8447 16507
rect 8389 16467 8447 16473
rect 8938 16464 8944 16516
rect 8996 16504 9002 16516
rect 12345 16507 12403 16513
rect 12345 16504 12357 16507
rect 8996 16476 12357 16504
rect 8996 16464 9002 16476
rect 12345 16473 12357 16476
rect 12391 16473 12403 16507
rect 12345 16467 12403 16473
rect 6920 16458 6972 16464
rect 4614 16396 4620 16448
rect 4672 16436 4678 16448
rect 4893 16439 4951 16445
rect 4893 16436 4905 16439
rect 4672 16408 4905 16436
rect 4672 16396 4678 16408
rect 4893 16405 4905 16408
rect 4939 16405 4951 16439
rect 4893 16399 4951 16405
rect 5169 16439 5227 16445
rect 5169 16405 5181 16439
rect 5215 16436 5227 16439
rect 5626 16436 5632 16448
rect 5215 16408 5632 16436
rect 5215 16405 5227 16408
rect 5169 16399 5227 16405
rect 5626 16396 5632 16408
rect 5684 16396 5690 16448
rect 7929 16439 7987 16445
rect 7929 16405 7941 16439
rect 7975 16436 7987 16439
rect 8478 16436 8484 16448
rect 7975 16408 8484 16436
rect 7975 16405 7987 16408
rect 7929 16399 7987 16405
rect 8478 16396 8484 16408
rect 8536 16396 8542 16448
rect 8754 16396 8760 16448
rect 8812 16396 8818 16448
rect 11146 16396 11152 16448
rect 11204 16436 11210 16448
rect 12452 16436 12480 16535
rect 12728 16504 12756 16535
rect 12894 16532 12900 16584
rect 12952 16532 12958 16584
rect 13262 16532 13268 16584
rect 13320 16532 13326 16584
rect 12728 16476 15424 16504
rect 11204 16408 12480 16436
rect 12621 16439 12679 16445
rect 11204 16396 11210 16408
rect 12621 16405 12633 16439
rect 12667 16436 12679 16439
rect 12802 16436 12808 16448
rect 12667 16408 12808 16436
rect 12667 16405 12679 16408
rect 12621 16399 12679 16405
rect 12802 16396 12808 16408
rect 12860 16396 12866 16448
rect 15396 16436 15424 16476
rect 15470 16464 15476 16516
rect 15528 16504 15534 16516
rect 17420 16504 17448 16612
rect 17512 16612 17632 16640
rect 17696 16680 18276 16708
rect 17512 16581 17540 16612
rect 17497 16575 17555 16581
rect 17497 16541 17509 16575
rect 17543 16541 17555 16575
rect 17497 16535 17555 16541
rect 17589 16575 17647 16581
rect 17589 16541 17601 16575
rect 17635 16572 17647 16575
rect 17696 16572 17724 16680
rect 18598 16668 18604 16720
rect 18656 16668 18662 16720
rect 19518 16708 19524 16720
rect 18800 16680 19524 16708
rect 17770 16600 17776 16652
rect 17828 16640 17834 16652
rect 17865 16643 17923 16649
rect 17865 16640 17877 16643
rect 17828 16612 17877 16640
rect 17828 16600 17834 16612
rect 17865 16609 17877 16612
rect 17911 16609 17923 16643
rect 18616 16640 18644 16668
rect 17865 16603 17923 16609
rect 18340 16612 18644 16640
rect 17635 16544 17724 16572
rect 17635 16541 17647 16544
rect 17589 16535 17647 16541
rect 17604 16504 17632 16535
rect 18046 16532 18052 16584
rect 18104 16532 18110 16584
rect 18340 16581 18368 16612
rect 18325 16575 18383 16581
rect 18325 16541 18337 16575
rect 18371 16541 18383 16575
rect 18325 16535 18383 16541
rect 18509 16575 18567 16581
rect 18509 16541 18521 16575
rect 18555 16541 18567 16575
rect 18509 16535 18567 16541
rect 18601 16575 18659 16581
rect 18601 16541 18613 16575
rect 18647 16541 18659 16575
rect 18601 16535 18659 16541
rect 18524 16504 18552 16535
rect 15528 16476 17382 16504
rect 17420 16476 17632 16504
rect 17977 16476 18552 16504
rect 18616 16504 18644 16535
rect 18690 16532 18696 16584
rect 18748 16532 18754 16584
rect 18800 16504 18828 16680
rect 19518 16668 19524 16680
rect 19576 16668 19582 16720
rect 20438 16668 20444 16720
rect 20496 16708 20502 16720
rect 20990 16708 20996 16720
rect 20496 16680 20996 16708
rect 20496 16668 20502 16680
rect 20990 16668 20996 16680
rect 21048 16668 21054 16720
rect 19242 16600 19248 16652
rect 19300 16640 19306 16652
rect 20530 16640 20536 16652
rect 19300 16612 20536 16640
rect 19300 16600 19306 16612
rect 20530 16600 20536 16612
rect 20588 16600 20594 16652
rect 20714 16600 20720 16652
rect 20772 16600 20778 16652
rect 21450 16640 21456 16652
rect 20916 16612 21456 16640
rect 18877 16575 18935 16581
rect 18877 16541 18889 16575
rect 18923 16572 18935 16575
rect 19058 16572 19064 16584
rect 18923 16544 19064 16572
rect 18923 16541 18935 16544
rect 18877 16535 18935 16541
rect 19058 16532 19064 16544
rect 19116 16532 19122 16584
rect 20438 16532 20444 16584
rect 20496 16532 20502 16584
rect 20548 16572 20576 16600
rect 20916 16572 20944 16612
rect 21284 16581 21312 16612
rect 21450 16600 21456 16612
rect 21508 16600 21514 16652
rect 25869 16643 25927 16649
rect 25869 16640 25881 16643
rect 22020 16612 25881 16640
rect 20548 16544 20944 16572
rect 20993 16575 21051 16581
rect 20993 16541 21005 16575
rect 21039 16541 21051 16575
rect 20993 16535 21051 16541
rect 21269 16575 21327 16581
rect 21269 16541 21281 16575
rect 21315 16541 21327 16575
rect 21269 16535 21327 16541
rect 21361 16575 21419 16581
rect 21361 16541 21373 16575
rect 21407 16541 21419 16575
rect 21361 16535 21419 16541
rect 21545 16575 21603 16581
rect 21545 16541 21557 16575
rect 21591 16572 21603 16575
rect 22020 16572 22048 16612
rect 21591 16544 22048 16572
rect 21591 16541 21603 16544
rect 21545 16535 21603 16541
rect 18616 16476 18828 16504
rect 20717 16507 20775 16513
rect 15528 16464 15534 16476
rect 16022 16436 16028 16448
rect 15396 16408 16028 16436
rect 16022 16396 16028 16408
rect 16080 16396 16086 16448
rect 17218 16396 17224 16448
rect 17276 16396 17282 16448
rect 17354 16436 17382 16476
rect 17977 16436 18005 16476
rect 17354 16408 18005 16436
rect 18046 16396 18052 16448
rect 18104 16396 18110 16448
rect 18524 16436 18552 16476
rect 20717 16473 20729 16507
rect 20763 16504 20775 16507
rect 21008 16504 21036 16535
rect 20763 16476 21036 16504
rect 20763 16473 20775 16476
rect 20717 16467 20775 16473
rect 21082 16464 21088 16516
rect 21140 16504 21146 16516
rect 21177 16507 21235 16513
rect 21177 16504 21189 16507
rect 21140 16476 21189 16504
rect 21140 16464 21146 16476
rect 21177 16473 21189 16476
rect 21223 16473 21235 16507
rect 21376 16504 21404 16535
rect 22094 16532 22100 16584
rect 22152 16532 22158 16584
rect 22204 16581 22232 16612
rect 25869 16609 25881 16612
rect 25915 16609 25927 16643
rect 25869 16603 25927 16609
rect 26142 16600 26148 16652
rect 26200 16600 26206 16652
rect 22189 16575 22247 16581
rect 22189 16541 22201 16575
rect 22235 16572 22247 16575
rect 23477 16575 23535 16581
rect 22235 16544 22269 16572
rect 22235 16541 22247 16544
rect 22189 16535 22247 16541
rect 23477 16541 23489 16575
rect 23523 16541 23535 16575
rect 23477 16535 23535 16541
rect 21177 16467 21235 16473
rect 21284 16476 21404 16504
rect 21284 16448 21312 16476
rect 21634 16464 21640 16516
rect 21692 16504 21698 16516
rect 23492 16504 23520 16535
rect 21692 16476 24440 16504
rect 21692 16464 21698 16476
rect 19702 16436 19708 16448
rect 18524 16408 19708 16436
rect 19702 16396 19708 16408
rect 19760 16396 19766 16448
rect 20809 16439 20867 16445
rect 20809 16405 20821 16439
rect 20855 16436 20867 16439
rect 20990 16436 20996 16448
rect 20855 16408 20996 16436
rect 20855 16405 20867 16408
rect 20809 16399 20867 16405
rect 20990 16396 20996 16408
rect 21048 16396 21054 16448
rect 21266 16396 21272 16448
rect 21324 16396 21330 16448
rect 21358 16396 21364 16448
rect 21416 16396 21422 16448
rect 23382 16396 23388 16448
rect 23440 16396 23446 16448
rect 24412 16445 24440 16476
rect 25314 16464 25320 16516
rect 25372 16464 25378 16516
rect 26602 16464 26608 16516
rect 26660 16464 26666 16516
rect 24397 16439 24455 16445
rect 24397 16405 24409 16439
rect 24443 16436 24455 16439
rect 24854 16436 24860 16448
rect 24443 16408 24860 16436
rect 24443 16405 24455 16408
rect 24397 16399 24455 16405
rect 24854 16396 24860 16408
rect 24912 16396 24918 16448
rect 1104 16346 28152 16368
rect 1104 16294 4874 16346
rect 4926 16294 4938 16346
rect 4990 16294 5002 16346
rect 5054 16294 5066 16346
rect 5118 16294 5130 16346
rect 5182 16294 28152 16346
rect 1104 16272 28152 16294
rect 6914 16232 6920 16244
rect 6748 16204 6920 16232
rect 1857 16099 1915 16105
rect 1857 16065 1869 16099
rect 1903 16096 1915 16099
rect 2498 16096 2504 16108
rect 1903 16068 2504 16096
rect 1903 16065 1915 16068
rect 1857 16059 1915 16065
rect 2498 16056 2504 16068
rect 2556 16056 2562 16108
rect 3878 16056 3884 16108
rect 3936 16056 3942 16108
rect 4614 16056 4620 16108
rect 4672 16056 4678 16108
rect 4890 16056 4896 16108
rect 4948 16056 4954 16108
rect 5350 16056 5356 16108
rect 5408 16056 5414 16108
rect 6748 16105 6776 16204
rect 6914 16192 6920 16204
rect 6972 16192 6978 16244
rect 16666 16232 16672 16244
rect 12406 16204 16672 16232
rect 8665 16167 8723 16173
rect 8665 16133 8677 16167
rect 8711 16164 8723 16167
rect 8754 16164 8760 16176
rect 8711 16136 8760 16164
rect 8711 16133 8723 16136
rect 8665 16127 8723 16133
rect 8754 16124 8760 16136
rect 8812 16124 8818 16176
rect 12406 16164 12434 16204
rect 16666 16192 16672 16204
rect 16724 16192 16730 16244
rect 16942 16192 16948 16244
rect 17000 16232 17006 16244
rect 17681 16235 17739 16241
rect 17681 16232 17693 16235
rect 17000 16204 17693 16232
rect 17000 16192 17006 16204
rect 17681 16201 17693 16204
rect 17727 16201 17739 16235
rect 17681 16195 17739 16201
rect 18506 16192 18512 16244
rect 18564 16232 18570 16244
rect 18782 16232 18788 16244
rect 18564 16204 18788 16232
rect 18564 16192 18570 16204
rect 18782 16192 18788 16204
rect 18840 16232 18846 16244
rect 19058 16232 19064 16244
rect 18840 16204 19064 16232
rect 18840 16192 18846 16204
rect 19058 16192 19064 16204
rect 19116 16232 19122 16244
rect 22002 16232 22008 16244
rect 19116 16204 22008 16232
rect 19116 16192 19122 16204
rect 22002 16192 22008 16204
rect 22060 16192 22066 16244
rect 22465 16235 22523 16241
rect 22465 16201 22477 16235
rect 22511 16232 22523 16235
rect 23477 16235 23535 16241
rect 23477 16232 23489 16235
rect 22511 16204 23489 16232
rect 22511 16201 22523 16204
rect 22465 16195 22523 16201
rect 23477 16201 23489 16204
rect 23523 16201 23535 16235
rect 23477 16195 23535 16201
rect 25314 16192 25320 16244
rect 25372 16232 25378 16244
rect 25682 16232 25688 16244
rect 25372 16204 25688 16232
rect 25372 16192 25378 16204
rect 25682 16192 25688 16204
rect 25740 16192 25746 16244
rect 9324 16136 9996 16164
rect 10902 16136 12434 16164
rect 6733 16099 6791 16105
rect 6733 16065 6745 16099
rect 6779 16065 6791 16099
rect 6733 16059 6791 16065
rect 7282 16056 7288 16108
rect 7340 16096 7346 16108
rect 7469 16099 7527 16105
rect 7469 16096 7481 16099
rect 7340 16068 7481 16096
rect 7340 16056 7346 16068
rect 7469 16065 7481 16068
rect 7515 16096 7527 16099
rect 8202 16096 8208 16108
rect 7515 16068 8208 16096
rect 7515 16065 7527 16068
rect 7469 16059 7527 16065
rect 8202 16056 8208 16068
rect 8260 16096 8266 16108
rect 8938 16096 8944 16108
rect 8260 16068 8944 16096
rect 8260 16056 8266 16068
rect 8938 16056 8944 16068
rect 8996 16056 9002 16108
rect 9030 16056 9036 16108
rect 9088 16056 9094 16108
rect 1949 16031 2007 16037
rect 1949 15997 1961 16031
rect 1995 16028 2007 16031
rect 2222 16028 2228 16040
rect 1995 16000 2228 16028
rect 1995 15997 2007 16000
rect 1949 15991 2007 15997
rect 2222 15988 2228 16000
rect 2280 15988 2286 16040
rect 4522 15988 4528 16040
rect 4580 15988 4586 16040
rect 8846 15988 8852 16040
rect 8904 15988 8910 16040
rect 9033 15963 9091 15969
rect 9033 15929 9045 15963
rect 9079 15960 9091 15963
rect 9324 15960 9352 16136
rect 9766 16056 9772 16108
rect 9824 16056 9830 16108
rect 9968 16105 9996 16136
rect 12802 16124 12808 16176
rect 12860 16124 12866 16176
rect 12986 16124 12992 16176
rect 13044 16124 13050 16176
rect 18141 16167 18199 16173
rect 18141 16133 18153 16167
rect 18187 16164 18199 16167
rect 18230 16164 18236 16176
rect 18187 16136 18236 16164
rect 18187 16133 18199 16136
rect 18141 16127 18199 16133
rect 18230 16124 18236 16136
rect 18288 16124 18294 16176
rect 18690 16124 18696 16176
rect 18748 16164 18754 16176
rect 22186 16164 22192 16176
rect 18748 16136 22192 16164
rect 18748 16124 18754 16136
rect 22186 16124 22192 16136
rect 22244 16124 22250 16176
rect 23382 16164 23388 16176
rect 23032 16136 23388 16164
rect 9953 16099 10011 16105
rect 9953 16065 9965 16099
rect 9999 16065 10011 16099
rect 13004 16096 13032 16124
rect 13081 16099 13139 16105
rect 13081 16096 13093 16099
rect 13004 16068 13093 16096
rect 9953 16059 10011 16065
rect 13081 16065 13093 16068
rect 13127 16065 13139 16099
rect 13081 16059 13139 16065
rect 17865 16099 17923 16105
rect 17865 16065 17877 16099
rect 17911 16096 17923 16099
rect 18046 16096 18052 16108
rect 17911 16068 18052 16096
rect 17911 16065 17923 16068
rect 17865 16059 17923 16065
rect 18046 16056 18052 16068
rect 18104 16056 18110 16108
rect 18506 16056 18512 16108
rect 18564 16056 18570 16108
rect 20530 16056 20536 16108
rect 20588 16056 20594 16108
rect 20806 16056 20812 16108
rect 20864 16056 20870 16108
rect 21266 16056 21272 16108
rect 21324 16056 21330 16108
rect 21453 16099 21511 16105
rect 21453 16065 21465 16099
rect 21499 16096 21511 16099
rect 21634 16096 21640 16108
rect 21499 16068 21640 16096
rect 21499 16065 21511 16068
rect 21453 16059 21511 16065
rect 21634 16056 21640 16068
rect 21692 16056 21698 16108
rect 22554 16096 22560 16108
rect 21744 16068 22560 16096
rect 12989 16031 13047 16037
rect 12989 15997 13001 16031
rect 13035 16028 13047 16031
rect 16850 16028 16856 16040
rect 13035 16000 16856 16028
rect 13035 15997 13047 16000
rect 12989 15991 13047 15997
rect 16850 15988 16856 16000
rect 16908 15988 16914 16040
rect 17954 15988 17960 16040
rect 18012 15988 18018 16040
rect 18233 16031 18291 16037
rect 18233 15997 18245 16031
rect 18279 16028 18291 16031
rect 18322 16028 18328 16040
rect 18279 16000 18328 16028
rect 18279 15997 18291 16000
rect 18233 15991 18291 15997
rect 18322 15988 18328 16000
rect 18380 15988 18386 16040
rect 20990 15988 20996 16040
rect 21048 16028 21054 16040
rect 21085 16031 21143 16037
rect 21085 16028 21097 16031
rect 21048 16000 21097 16028
rect 21048 15988 21054 16000
rect 21085 15997 21097 16000
rect 21131 15997 21143 16031
rect 21085 15991 21143 15997
rect 9079 15932 9352 15960
rect 13265 15963 13323 15969
rect 9079 15929 9091 15932
rect 9033 15923 9091 15929
rect 13265 15929 13277 15963
rect 13311 15960 13323 15963
rect 17034 15960 17040 15972
rect 13311 15932 17040 15960
rect 13311 15929 13323 15932
rect 13265 15923 13323 15929
rect 17034 15920 17040 15932
rect 17092 15920 17098 15972
rect 17402 15920 17408 15972
rect 17460 15960 17466 15972
rect 18417 15963 18475 15969
rect 18417 15960 18429 15963
rect 17460 15932 18429 15960
rect 17460 15920 17466 15932
rect 18417 15929 18429 15932
rect 18463 15929 18475 15963
rect 18417 15923 18475 15929
rect 18690 15920 18696 15972
rect 18748 15960 18754 15972
rect 21744 15960 21772 16068
rect 22554 16056 22560 16068
rect 22612 16096 22618 16108
rect 22649 16099 22707 16105
rect 22649 16096 22661 16099
rect 22612 16068 22661 16096
rect 22612 16056 22618 16068
rect 22649 16065 22661 16068
rect 22695 16065 22707 16099
rect 22649 16059 22707 16065
rect 22738 16056 22744 16108
rect 22796 16056 22802 16108
rect 22922 16056 22928 16108
rect 22980 16056 22986 16108
rect 23032 16105 23060 16136
rect 23382 16124 23388 16136
rect 23440 16164 23446 16176
rect 23753 16167 23811 16173
rect 23753 16164 23765 16167
rect 23440 16136 23765 16164
rect 23440 16124 23446 16136
rect 23753 16133 23765 16136
rect 23799 16133 23811 16167
rect 23753 16127 23811 16133
rect 25498 16124 25504 16176
rect 25556 16164 25562 16176
rect 25593 16167 25651 16173
rect 25593 16164 25605 16167
rect 25556 16136 25605 16164
rect 25556 16124 25562 16136
rect 25593 16133 25605 16136
rect 25639 16133 25651 16167
rect 25593 16127 25651 16133
rect 23017 16099 23075 16105
rect 23017 16065 23029 16099
rect 23063 16065 23075 16099
rect 23017 16059 23075 16065
rect 23293 16099 23351 16105
rect 23293 16065 23305 16099
rect 23339 16065 23351 16099
rect 23293 16059 23351 16065
rect 22094 15988 22100 16040
rect 22152 16028 22158 16040
rect 23109 16031 23167 16037
rect 23109 16028 23121 16031
rect 22152 16000 23121 16028
rect 22152 15988 22158 16000
rect 23109 15997 23121 16000
rect 23155 15997 23167 16031
rect 23109 15991 23167 15997
rect 18748 15932 21772 15960
rect 18748 15920 18754 15932
rect 2133 15895 2191 15901
rect 2133 15861 2145 15895
rect 2179 15892 2191 15895
rect 2314 15892 2320 15904
rect 2179 15864 2320 15892
rect 2179 15861 2191 15864
rect 2133 15855 2191 15861
rect 2314 15852 2320 15864
rect 2372 15852 2378 15904
rect 8205 15895 8263 15901
rect 8205 15861 8217 15895
rect 8251 15892 8263 15895
rect 8294 15892 8300 15904
rect 8251 15864 8300 15892
rect 8251 15861 8263 15864
rect 8205 15855 8263 15861
rect 8294 15852 8300 15864
rect 8352 15852 8358 15904
rect 12802 15852 12808 15904
rect 12860 15852 12866 15904
rect 18138 15852 18144 15904
rect 18196 15852 18202 15904
rect 18509 15895 18567 15901
rect 18509 15861 18521 15895
rect 18555 15892 18567 15895
rect 18598 15892 18604 15904
rect 18555 15864 18604 15892
rect 18555 15861 18567 15864
rect 18509 15855 18567 15861
rect 18598 15852 18604 15864
rect 18656 15852 18662 15904
rect 19245 15895 19303 15901
rect 19245 15861 19257 15895
rect 19291 15892 19303 15895
rect 19334 15892 19340 15904
rect 19291 15864 19340 15892
rect 19291 15861 19303 15864
rect 19245 15855 19303 15861
rect 19334 15852 19340 15864
rect 19392 15852 19398 15904
rect 19794 15852 19800 15904
rect 19852 15892 19858 15904
rect 20625 15895 20683 15901
rect 20625 15892 20637 15895
rect 19852 15864 20637 15892
rect 19852 15852 19858 15864
rect 20625 15861 20637 15864
rect 20671 15861 20683 15895
rect 20625 15855 20683 15861
rect 20993 15895 21051 15901
rect 20993 15861 21005 15895
rect 21039 15892 21051 15895
rect 21082 15892 21088 15904
rect 21039 15864 21088 15892
rect 21039 15861 21051 15864
rect 20993 15855 21051 15861
rect 21082 15852 21088 15864
rect 21140 15852 21146 15904
rect 21269 15895 21327 15901
rect 21269 15861 21281 15895
rect 21315 15892 21327 15895
rect 21358 15892 21364 15904
rect 21315 15864 21364 15892
rect 21315 15861 21327 15864
rect 21269 15855 21327 15861
rect 21358 15852 21364 15864
rect 21416 15852 21422 15904
rect 23308 15892 23336 16059
rect 23566 16056 23572 16108
rect 23624 16056 23630 16108
rect 23661 16099 23719 16105
rect 23661 16065 23673 16099
rect 23707 16065 23719 16099
rect 23661 16059 23719 16065
rect 23382 15988 23388 16040
rect 23440 16028 23446 16040
rect 23676 16028 23704 16059
rect 23842 16056 23848 16108
rect 23900 16096 23906 16108
rect 23937 16099 23995 16105
rect 23937 16096 23949 16099
rect 23900 16068 23949 16096
rect 23900 16056 23906 16068
rect 23937 16065 23949 16068
rect 23983 16065 23995 16099
rect 23937 16059 23995 16065
rect 23440 16000 23704 16028
rect 23440 15988 23446 16000
rect 24121 15895 24179 15901
rect 24121 15892 24133 15895
rect 23308 15864 24133 15892
rect 24121 15861 24133 15864
rect 24167 15861 24179 15895
rect 24121 15855 24179 15861
rect 1104 15802 28152 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 28152 15802
rect 1104 15728 28152 15750
rect 7558 15648 7564 15700
rect 7616 15648 7622 15700
rect 16942 15648 16948 15700
rect 17000 15688 17006 15700
rect 18690 15688 18696 15700
rect 17000 15660 18696 15688
rect 17000 15648 17006 15660
rect 18690 15648 18696 15660
rect 18748 15648 18754 15700
rect 20901 15691 20959 15697
rect 20901 15657 20913 15691
rect 20947 15657 20959 15691
rect 20901 15651 20959 15657
rect 8478 15620 8484 15632
rect 7760 15592 8484 15620
rect 4525 15555 4583 15561
rect 4525 15521 4537 15555
rect 4571 15552 4583 15555
rect 4614 15552 4620 15564
rect 4571 15524 4620 15552
rect 4571 15521 4583 15524
rect 4525 15515 4583 15521
rect 4614 15512 4620 15524
rect 4672 15512 4678 15564
rect 1394 15444 1400 15496
rect 1452 15444 1458 15496
rect 2774 15444 2780 15496
rect 2832 15444 2838 15496
rect 3053 15487 3111 15493
rect 3053 15453 3065 15487
rect 3099 15484 3111 15487
rect 3234 15484 3240 15496
rect 3099 15456 3240 15484
rect 3099 15453 3111 15456
rect 3053 15447 3111 15453
rect 3234 15444 3240 15456
rect 3292 15444 3298 15496
rect 4433 15487 4491 15493
rect 4433 15453 4445 15487
rect 4479 15453 4491 15487
rect 4433 15447 4491 15453
rect 1673 15419 1731 15425
rect 1673 15385 1685 15419
rect 1719 15416 1731 15419
rect 2038 15416 2044 15428
rect 1719 15388 2044 15416
rect 1719 15385 1731 15388
rect 1673 15379 1731 15385
rect 2038 15376 2044 15388
rect 2096 15376 2102 15428
rect 4448 15416 4476 15447
rect 4890 15444 4896 15496
rect 4948 15444 4954 15496
rect 5077 15487 5135 15493
rect 5077 15453 5089 15487
rect 5123 15484 5135 15487
rect 5350 15484 5356 15496
rect 5123 15456 5356 15484
rect 5123 15453 5135 15456
rect 5077 15447 5135 15453
rect 5350 15444 5356 15456
rect 5408 15444 5414 15496
rect 7760 15493 7788 15592
rect 8478 15580 8484 15592
rect 8536 15580 8542 15632
rect 8665 15623 8723 15629
rect 8665 15589 8677 15623
rect 8711 15620 8723 15623
rect 8846 15620 8852 15632
rect 8711 15592 8852 15620
rect 8711 15589 8723 15592
rect 8665 15583 8723 15589
rect 8846 15580 8852 15592
rect 8904 15580 8910 15632
rect 19426 15580 19432 15632
rect 19484 15580 19490 15632
rect 20349 15623 20407 15629
rect 20349 15620 20361 15623
rect 19628 15592 20361 15620
rect 8021 15555 8079 15561
rect 8021 15521 8033 15555
rect 8067 15552 8079 15555
rect 8294 15552 8300 15564
rect 8067 15524 8300 15552
rect 8067 15521 8079 15524
rect 8021 15515 8079 15521
rect 8294 15512 8300 15524
rect 8352 15512 8358 15564
rect 7745 15487 7803 15493
rect 7745 15453 7757 15487
rect 7791 15453 7803 15487
rect 7745 15447 7803 15453
rect 7837 15487 7895 15493
rect 7837 15453 7849 15487
rect 7883 15484 7895 15487
rect 7926 15484 7932 15496
rect 7883 15456 7932 15484
rect 7883 15453 7895 15456
rect 7837 15447 7895 15453
rect 7926 15444 7932 15456
rect 7984 15444 7990 15496
rect 8113 15487 8171 15493
rect 8113 15453 8125 15487
rect 8159 15484 8171 15487
rect 8386 15484 8392 15496
rect 8159 15456 8392 15484
rect 8159 15453 8171 15456
rect 8113 15447 8171 15453
rect 8386 15444 8392 15456
rect 8444 15444 8450 15496
rect 8570 15444 8576 15496
rect 8628 15444 8634 15496
rect 8754 15444 8760 15496
rect 8812 15444 8818 15496
rect 8864 15484 8892 15580
rect 19628 15564 19656 15592
rect 20349 15589 20361 15592
rect 20395 15589 20407 15623
rect 20916 15620 20944 15651
rect 21082 15648 21088 15700
rect 21140 15648 21146 15700
rect 21266 15648 21272 15700
rect 21324 15688 21330 15700
rect 23477 15691 23535 15697
rect 21324 15660 21956 15688
rect 21324 15648 21330 15660
rect 21358 15620 21364 15632
rect 20916 15592 21364 15620
rect 20349 15583 20407 15589
rect 21358 15580 21364 15592
rect 21416 15580 21422 15632
rect 9030 15512 9036 15564
rect 9088 15552 9094 15564
rect 9088 15524 9444 15552
rect 9088 15512 9094 15524
rect 9309 15487 9367 15493
rect 9309 15484 9321 15487
rect 8864 15456 9321 15484
rect 9309 15453 9321 15456
rect 9355 15453 9367 15487
rect 9416 15484 9444 15524
rect 19610 15512 19616 15564
rect 19668 15512 19674 15564
rect 20990 15552 20996 15564
rect 20548 15524 20996 15552
rect 9858 15484 9864 15496
rect 9416 15456 9864 15484
rect 9309 15447 9367 15453
rect 9858 15444 9864 15456
rect 9916 15444 9922 15496
rect 19426 15444 19432 15496
rect 19484 15444 19490 15496
rect 19794 15444 19800 15496
rect 19852 15444 19858 15496
rect 20548 15493 20576 15524
rect 20990 15512 20996 15524
rect 21048 15512 21054 15564
rect 21100 15524 21496 15552
rect 20533 15487 20591 15493
rect 20533 15453 20545 15487
rect 20579 15453 20591 15487
rect 20533 15447 20591 15453
rect 20714 15444 20720 15496
rect 20772 15444 20778 15496
rect 21100 15484 21128 15524
rect 21468 15496 21496 15524
rect 20916 15456 21128 15484
rect 4985 15419 5043 15425
rect 4985 15416 4997 15419
rect 4448 15388 4997 15416
rect 4985 15385 4997 15388
rect 5031 15385 5043 15419
rect 8588 15416 8616 15444
rect 9122 15416 9128 15428
rect 8588 15388 9128 15416
rect 4985 15379 5043 15385
rect 9122 15376 9128 15388
rect 9180 15376 9186 15428
rect 20916 15416 20944 15456
rect 21266 15444 21272 15496
rect 21324 15444 21330 15496
rect 21450 15444 21456 15496
rect 21508 15444 21514 15496
rect 21545 15487 21603 15493
rect 21545 15453 21557 15487
rect 21591 15453 21603 15487
rect 21545 15447 21603 15453
rect 10810 15388 20944 15416
rect 20993 15419 21051 15425
rect 20993 15385 21005 15419
rect 21039 15416 21051 15419
rect 21560 15416 21588 15447
rect 21634 15444 21640 15496
rect 21692 15484 21698 15496
rect 21928 15493 21956 15660
rect 23477 15657 23489 15691
rect 23523 15688 23535 15691
rect 23566 15688 23572 15700
rect 23523 15660 23572 15688
rect 23523 15657 23535 15660
rect 23477 15651 23535 15657
rect 23566 15648 23572 15660
rect 23624 15648 23630 15700
rect 23937 15691 23995 15697
rect 23937 15657 23949 15691
rect 23983 15688 23995 15691
rect 24397 15691 24455 15697
rect 24397 15688 24409 15691
rect 23983 15660 24409 15688
rect 23983 15657 23995 15660
rect 23937 15651 23995 15657
rect 24397 15657 24409 15660
rect 24443 15688 24455 15691
rect 24486 15688 24492 15700
rect 24443 15660 24492 15688
rect 24443 15657 24455 15660
rect 24397 15651 24455 15657
rect 24486 15648 24492 15660
rect 24544 15648 24550 15700
rect 24578 15648 24584 15700
rect 24636 15648 24642 15700
rect 22370 15580 22376 15632
rect 22428 15620 22434 15632
rect 22646 15620 22652 15632
rect 22428 15592 22652 15620
rect 22428 15580 22434 15592
rect 22646 15580 22652 15592
rect 22704 15620 22710 15632
rect 22922 15620 22928 15632
rect 22704 15592 22928 15620
rect 22704 15580 22710 15592
rect 22922 15580 22928 15592
rect 22980 15620 22986 15632
rect 23109 15623 23167 15629
rect 23109 15620 23121 15623
rect 22980 15592 23121 15620
rect 22980 15580 22986 15592
rect 23109 15589 23121 15592
rect 23155 15589 23167 15623
rect 23109 15583 23167 15589
rect 23845 15623 23903 15629
rect 23845 15589 23857 15623
rect 23891 15620 23903 15623
rect 24857 15623 24915 15629
rect 24857 15620 24869 15623
rect 23891 15592 24869 15620
rect 23891 15589 23903 15592
rect 23845 15583 23903 15589
rect 24857 15589 24869 15592
rect 24903 15589 24915 15623
rect 24857 15583 24915 15589
rect 24578 15512 24584 15564
rect 24636 15552 24642 15564
rect 24636 15524 25084 15552
rect 24636 15512 24642 15524
rect 21729 15487 21787 15493
rect 21729 15484 21741 15487
rect 21692 15456 21741 15484
rect 21692 15444 21698 15456
rect 21729 15453 21741 15456
rect 21775 15453 21787 15487
rect 21729 15447 21787 15453
rect 21913 15487 21971 15493
rect 21913 15453 21925 15487
rect 21959 15484 21971 15487
rect 22094 15484 22100 15496
rect 21959 15456 22100 15484
rect 21959 15453 21971 15456
rect 21913 15447 21971 15453
rect 22094 15444 22100 15456
rect 22152 15444 22158 15496
rect 22925 15487 22983 15493
rect 22925 15453 22937 15487
rect 22971 15453 22983 15487
rect 22925 15447 22983 15453
rect 21821 15419 21879 15425
rect 21821 15416 21833 15419
rect 21039 15388 21833 15416
rect 21039 15385 21051 15388
rect 20993 15379 21051 15385
rect 21821 15385 21833 15388
rect 21867 15385 21879 15419
rect 21821 15379 21879 15385
rect 3234 15308 3240 15360
rect 3292 15348 3298 15360
rect 3421 15351 3479 15357
rect 3421 15348 3433 15351
rect 3292 15320 3433 15348
rect 3292 15308 3298 15320
rect 3421 15317 3433 15320
rect 3467 15317 3479 15351
rect 3421 15311 3479 15317
rect 4798 15308 4804 15360
rect 4856 15308 4862 15360
rect 18598 15308 18604 15360
rect 18656 15348 18662 15360
rect 22940 15348 22968 15447
rect 23198 15444 23204 15496
rect 23256 15484 23262 15496
rect 23750 15484 23756 15496
rect 23256 15456 23756 15484
rect 23256 15444 23262 15456
rect 23750 15444 23756 15456
rect 23808 15444 23814 15496
rect 24026 15444 24032 15496
rect 24084 15444 24090 15496
rect 24210 15444 24216 15496
rect 24268 15444 24274 15496
rect 25056 15493 25084 15524
rect 25041 15487 25099 15493
rect 24596 15456 24992 15484
rect 24596 15357 24624 15456
rect 24765 15419 24823 15425
rect 24765 15385 24777 15419
rect 24811 15416 24823 15419
rect 24854 15416 24860 15428
rect 24811 15388 24860 15416
rect 24811 15385 24823 15388
rect 24765 15379 24823 15385
rect 24854 15376 24860 15388
rect 24912 15376 24918 15428
rect 24964 15416 24992 15456
rect 25041 15453 25053 15487
rect 25087 15453 25099 15487
rect 25041 15447 25099 15453
rect 25130 15444 25136 15496
rect 25188 15444 25194 15496
rect 25148 15416 25176 15444
rect 24964 15388 25176 15416
rect 18656 15320 22968 15348
rect 24565 15351 24624 15357
rect 18656 15308 18662 15320
rect 24565 15317 24577 15351
rect 24611 15320 24624 15351
rect 24611 15317 24623 15320
rect 24565 15311 24623 15317
rect 1104 15258 28152 15280
rect 1104 15206 4874 15258
rect 4926 15206 4938 15258
rect 4990 15206 5002 15258
rect 5054 15206 5066 15258
rect 5118 15206 5130 15258
rect 5182 15206 28152 15258
rect 1104 15184 28152 15206
rect 2774 15104 2780 15156
rect 2832 15144 2838 15156
rect 2869 15147 2927 15153
rect 2869 15144 2881 15147
rect 2832 15116 2881 15144
rect 2832 15104 2838 15116
rect 2869 15113 2881 15116
rect 2915 15113 2927 15147
rect 2869 15107 2927 15113
rect 12069 15147 12127 15153
rect 12069 15113 12081 15147
rect 12115 15144 12127 15147
rect 12802 15144 12808 15156
rect 12115 15116 12808 15144
rect 12115 15113 12127 15116
rect 12069 15107 12127 15113
rect 12802 15104 12808 15116
rect 12860 15104 12866 15156
rect 14826 15104 14832 15156
rect 14884 15144 14890 15156
rect 15105 15147 15163 15153
rect 15105 15144 15117 15147
rect 14884 15116 15117 15144
rect 14884 15104 14890 15116
rect 15105 15113 15117 15116
rect 15151 15113 15163 15147
rect 15105 15107 15163 15113
rect 18506 15104 18512 15156
rect 18564 15144 18570 15156
rect 18877 15147 18935 15153
rect 18877 15144 18889 15147
rect 18564 15116 18889 15144
rect 18564 15104 18570 15116
rect 18877 15113 18889 15116
rect 18923 15113 18935 15147
rect 18877 15107 18935 15113
rect 20714 15104 20720 15156
rect 20772 15144 20778 15156
rect 20809 15147 20867 15153
rect 20809 15144 20821 15147
rect 20772 15116 20821 15144
rect 20772 15104 20778 15116
rect 20809 15113 20821 15116
rect 20855 15113 20867 15147
rect 20809 15107 20867 15113
rect 5350 15076 5356 15088
rect 2976 15048 5356 15076
rect 2976 15017 3004 15048
rect 5350 15036 5356 15048
rect 5408 15036 5414 15088
rect 9858 15036 9864 15088
rect 9916 15036 9922 15088
rect 10226 15036 10232 15088
rect 10284 15076 10290 15088
rect 11793 15079 11851 15085
rect 11793 15076 11805 15079
rect 10284 15048 11805 15076
rect 10284 15036 10290 15048
rect 11793 15045 11805 15048
rect 11839 15045 11851 15079
rect 11793 15039 11851 15045
rect 15289 15079 15347 15085
rect 15289 15045 15301 15079
rect 15335 15076 15347 15079
rect 22002 15076 22008 15088
rect 15335 15048 22008 15076
rect 15335 15045 15347 15048
rect 15289 15039 15347 15045
rect 22002 15036 22008 15048
rect 22060 15036 22066 15088
rect 2777 15011 2835 15017
rect 2777 14977 2789 15011
rect 2823 14977 2835 15011
rect 2777 14971 2835 14977
rect 2961 15011 3019 15017
rect 2961 14977 2973 15011
rect 3007 14977 3019 15011
rect 2961 14971 3019 14977
rect 2038 14900 2044 14952
rect 2096 14940 2102 14952
rect 2792 14940 2820 14971
rect 3142 14968 3148 15020
rect 3200 15008 3206 15020
rect 3237 15011 3295 15017
rect 3237 15008 3249 15011
rect 3200 14980 3249 15008
rect 3200 14968 3206 14980
rect 3237 14977 3249 14980
rect 3283 15008 3295 15011
rect 7650 15008 7656 15020
rect 3283 14980 7656 15008
rect 3283 14977 3295 14980
rect 3237 14971 3295 14977
rect 7650 14968 7656 14980
rect 7708 14968 7714 15020
rect 8205 15011 8263 15017
rect 8205 14977 8217 15011
rect 8251 15008 8263 15011
rect 8294 15008 8300 15020
rect 8251 14980 8300 15008
rect 8251 14977 8263 14980
rect 8205 14971 8263 14977
rect 8294 14968 8300 14980
rect 8352 14968 8358 15020
rect 8386 14968 8392 15020
rect 8444 14968 8450 15020
rect 11514 14968 11520 15020
rect 11572 14968 11578 15020
rect 11698 14968 11704 15020
rect 11756 14968 11762 15020
rect 11882 14968 11888 15020
rect 11940 14968 11946 15020
rect 12618 14968 12624 15020
rect 12676 14968 12682 15020
rect 12989 15011 13047 15017
rect 12989 14977 13001 15011
rect 13035 15008 13047 15011
rect 13630 15008 13636 15020
rect 13035 14980 13636 15008
rect 13035 14977 13047 14980
rect 12989 14971 13047 14977
rect 13630 14968 13636 14980
rect 13688 14968 13694 15020
rect 14274 14968 14280 15020
rect 14332 15008 14338 15020
rect 14332 14980 15700 15008
rect 14332 14968 14338 14980
rect 3160 14940 3188 14968
rect 2096 14912 3188 14940
rect 2096 14900 2102 14912
rect 5442 14900 5448 14952
rect 5500 14900 5506 14952
rect 12161 14943 12219 14949
rect 12161 14909 12173 14943
rect 12207 14909 12219 14943
rect 12161 14903 12219 14909
rect 12713 14943 12771 14949
rect 12713 14909 12725 14943
rect 12759 14909 12771 14943
rect 12713 14903 12771 14909
rect 12897 14943 12955 14949
rect 12897 14909 12909 14943
rect 12943 14940 12955 14943
rect 13170 14940 13176 14952
rect 12943 14912 13176 14940
rect 12943 14909 12955 14912
rect 12897 14903 12955 14909
rect 4798 14832 4804 14884
rect 4856 14872 4862 14884
rect 5721 14875 5779 14881
rect 5721 14872 5733 14875
rect 4856 14844 5733 14872
rect 4856 14832 4862 14844
rect 5721 14841 5733 14844
rect 5767 14841 5779 14875
rect 5721 14835 5779 14841
rect 3142 14764 3148 14816
rect 3200 14804 3206 14816
rect 3329 14807 3387 14813
rect 3329 14804 3341 14807
rect 3200 14776 3341 14804
rect 3200 14764 3206 14776
rect 3329 14773 3341 14776
rect 3375 14804 3387 14807
rect 4614 14804 4620 14816
rect 3375 14776 4620 14804
rect 3375 14773 3387 14776
rect 3329 14767 3387 14773
rect 4614 14764 4620 14776
rect 4672 14764 4678 14816
rect 5905 14807 5963 14813
rect 5905 14773 5917 14807
rect 5951 14804 5963 14807
rect 6178 14804 6184 14816
rect 5951 14776 6184 14804
rect 5951 14773 5963 14776
rect 5905 14767 5963 14773
rect 6178 14764 6184 14776
rect 6236 14764 6242 14816
rect 12176 14804 12204 14903
rect 12250 14832 12256 14884
rect 12308 14832 12314 14884
rect 12728 14872 12756 14903
rect 13170 14900 13176 14912
rect 13228 14940 13234 14952
rect 13998 14940 14004 14952
rect 13228 14912 14004 14940
rect 13228 14900 13234 14912
rect 13998 14900 14004 14912
rect 14056 14900 14062 14952
rect 15194 14900 15200 14952
rect 15252 14900 15258 14952
rect 15286 14900 15292 14952
rect 15344 14940 15350 14952
rect 15672 14949 15700 14980
rect 18138 14968 18144 15020
rect 18196 15008 18202 15020
rect 18417 15011 18475 15017
rect 18417 15008 18429 15011
rect 18196 14980 18429 15008
rect 18196 14968 18202 14980
rect 18417 14977 18429 14980
rect 18463 14977 18475 15011
rect 18417 14971 18475 14977
rect 18693 15011 18751 15017
rect 18693 14977 18705 15011
rect 18739 15008 18751 15011
rect 19610 15008 19616 15020
rect 18739 14980 19616 15008
rect 18739 14977 18751 14980
rect 18693 14971 18751 14977
rect 19610 14968 19616 14980
rect 19668 14968 19674 15020
rect 21177 15011 21235 15017
rect 21177 14977 21189 15011
rect 21223 15008 21235 15011
rect 21266 15008 21272 15020
rect 21223 14980 21272 15008
rect 21223 14977 21235 14980
rect 21177 14971 21235 14977
rect 21266 14968 21272 14980
rect 21324 15008 21330 15020
rect 24305 15011 24363 15017
rect 21324 14980 23060 15008
rect 21324 14968 21330 14980
rect 15381 14943 15439 14949
rect 15381 14940 15393 14943
rect 15344 14912 15393 14940
rect 15344 14900 15350 14912
rect 15381 14909 15393 14912
rect 15427 14909 15439 14943
rect 15381 14903 15439 14909
rect 15657 14943 15715 14949
rect 15657 14909 15669 14943
rect 15703 14940 15715 14943
rect 16850 14940 16856 14952
rect 15703 14912 16856 14940
rect 15703 14909 15715 14912
rect 15657 14903 15715 14909
rect 16850 14900 16856 14912
rect 16908 14900 16914 14952
rect 18322 14900 18328 14952
rect 18380 14940 18386 14952
rect 18509 14943 18567 14949
rect 18509 14940 18521 14943
rect 18380 14912 18521 14940
rect 18380 14900 18386 14912
rect 18509 14909 18521 14912
rect 18555 14909 18567 14943
rect 18509 14903 18567 14909
rect 21085 14943 21143 14949
rect 21085 14909 21097 14943
rect 21131 14940 21143 14943
rect 21450 14940 21456 14952
rect 21131 14912 21456 14940
rect 21131 14909 21143 14912
rect 21085 14903 21143 14909
rect 21450 14900 21456 14912
rect 21508 14940 21514 14952
rect 21818 14940 21824 14952
rect 21508 14912 21824 14940
rect 21508 14900 21514 14912
rect 21818 14900 21824 14912
rect 21876 14900 21882 14952
rect 13446 14872 13452 14884
rect 12728 14844 13452 14872
rect 13446 14832 13452 14844
rect 13504 14832 13510 14884
rect 23032 14816 23060 14980
rect 24305 14977 24317 15011
rect 24351 15008 24363 15011
rect 24578 15008 24584 15020
rect 24351 14980 24584 15008
rect 24351 14977 24363 14980
rect 24305 14971 24363 14977
rect 24578 14968 24584 14980
rect 24636 14968 24642 15020
rect 14182 14804 14188 14816
rect 12176 14776 14188 14804
rect 14182 14764 14188 14776
rect 14240 14764 14246 14816
rect 15562 14764 15568 14816
rect 15620 14804 15626 14816
rect 15930 14804 15936 14816
rect 15620 14776 15936 14804
rect 15620 14764 15626 14776
rect 15930 14764 15936 14776
rect 15988 14764 15994 14816
rect 18693 14807 18751 14813
rect 18693 14773 18705 14807
rect 18739 14804 18751 14807
rect 20070 14804 20076 14816
rect 18739 14776 20076 14804
rect 18739 14773 18751 14776
rect 18693 14767 18751 14773
rect 20070 14764 20076 14776
rect 20128 14764 20134 14816
rect 23014 14764 23020 14816
rect 23072 14804 23078 14816
rect 24213 14807 24271 14813
rect 24213 14804 24225 14807
rect 23072 14776 24225 14804
rect 23072 14764 23078 14776
rect 24213 14773 24225 14776
rect 24259 14773 24271 14807
rect 24213 14767 24271 14773
rect 1104 14714 28152 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 28152 14714
rect 1104 14640 28152 14662
rect 11974 14560 11980 14612
rect 12032 14600 12038 14612
rect 12032 14572 12572 14600
rect 12032 14560 12038 14572
rect 3973 14535 4031 14541
rect 3973 14532 3985 14535
rect 3528 14504 3985 14532
rect 3528 14473 3556 14504
rect 3973 14501 3985 14504
rect 4019 14532 4031 14535
rect 4706 14532 4712 14544
rect 4019 14504 4712 14532
rect 4019 14501 4031 14504
rect 3973 14495 4031 14501
rect 4706 14492 4712 14504
rect 4764 14492 4770 14544
rect 6457 14535 6515 14541
rect 6457 14501 6469 14535
rect 6503 14532 6515 14535
rect 8386 14532 8392 14544
rect 6503 14504 8392 14532
rect 6503 14501 6515 14504
rect 6457 14495 6515 14501
rect 8386 14492 8392 14504
rect 8444 14492 8450 14544
rect 12544 14532 12572 14572
rect 12618 14560 12624 14612
rect 12676 14600 12682 14612
rect 13081 14603 13139 14609
rect 13081 14600 13093 14603
rect 12676 14572 13093 14600
rect 12676 14560 12682 14572
rect 13081 14569 13093 14572
rect 13127 14569 13139 14603
rect 13081 14563 13139 14569
rect 14182 14560 14188 14612
rect 14240 14600 14246 14612
rect 15102 14600 15108 14612
rect 14240 14572 15108 14600
rect 14240 14560 14246 14572
rect 15102 14560 15108 14572
rect 15160 14600 15166 14612
rect 15565 14603 15623 14609
rect 15160 14572 15516 14600
rect 15160 14560 15166 14572
rect 14691 14535 14749 14541
rect 14691 14532 14703 14535
rect 12544 14504 13400 14532
rect 3513 14467 3571 14473
rect 3513 14433 3525 14467
rect 3559 14433 3571 14467
rect 3513 14427 3571 14433
rect 4065 14467 4123 14473
rect 4065 14433 4077 14467
rect 4111 14464 4123 14467
rect 4246 14464 4252 14476
rect 4111 14436 4252 14464
rect 4111 14433 4123 14436
rect 4065 14427 4123 14433
rect 4246 14424 4252 14436
rect 4304 14424 4310 14476
rect 4341 14467 4399 14473
rect 4341 14433 4353 14467
rect 4387 14464 4399 14467
rect 4387 14436 5488 14464
rect 4387 14433 4399 14436
rect 4341 14427 4399 14433
rect 5460 14408 5488 14436
rect 5902 14424 5908 14476
rect 5960 14464 5966 14476
rect 6089 14467 6147 14473
rect 6089 14464 6101 14467
rect 5960 14436 6101 14464
rect 5960 14424 5966 14436
rect 6089 14433 6101 14436
rect 6135 14464 6147 14467
rect 7009 14467 7067 14473
rect 7009 14464 7021 14467
rect 6135 14436 7021 14464
rect 6135 14433 6147 14436
rect 6089 14427 6147 14433
rect 7009 14433 7021 14436
rect 7055 14433 7067 14467
rect 7009 14427 7067 14433
rect 11057 14467 11115 14473
rect 11057 14433 11069 14467
rect 11103 14464 11115 14467
rect 11882 14464 11888 14476
rect 11103 14436 11888 14464
rect 11103 14433 11115 14436
rect 11057 14427 11115 14433
rect 11882 14424 11888 14436
rect 11940 14424 11946 14476
rect 12710 14424 12716 14476
rect 12768 14464 12774 14476
rect 12768 14436 13308 14464
rect 12768 14424 12774 14436
rect 2774 14356 2780 14408
rect 2832 14356 2838 14408
rect 3234 14356 3240 14408
rect 3292 14356 3298 14408
rect 3602 14356 3608 14408
rect 3660 14396 3666 14408
rect 3881 14399 3939 14405
rect 3881 14396 3893 14399
rect 3660 14368 3893 14396
rect 3660 14356 3666 14368
rect 3881 14365 3893 14368
rect 3927 14365 3939 14399
rect 3881 14359 3939 14365
rect 4154 14356 4160 14408
rect 4212 14396 4218 14408
rect 4614 14396 4620 14408
rect 4212 14368 4620 14396
rect 4212 14356 4218 14368
rect 4614 14356 4620 14368
rect 4672 14356 4678 14408
rect 4798 14356 4804 14408
rect 4856 14396 4862 14408
rect 5077 14399 5135 14405
rect 5077 14396 5089 14399
rect 4856 14368 5089 14396
rect 4856 14356 4862 14368
rect 5077 14365 5089 14368
rect 5123 14365 5135 14399
rect 5077 14359 5135 14365
rect 5442 14356 5448 14408
rect 5500 14356 5506 14408
rect 6178 14356 6184 14408
rect 6236 14356 6242 14408
rect 6730 14356 6736 14408
rect 6788 14356 6794 14408
rect 11146 14356 11152 14408
rect 11204 14356 11210 14408
rect 11238 14356 11244 14408
rect 11296 14356 11302 14408
rect 13280 14405 13308 14436
rect 13372 14405 13400 14504
rect 14292 14504 14703 14532
rect 13817 14467 13875 14473
rect 13817 14464 13829 14467
rect 13648 14436 13829 14464
rect 13648 14408 13676 14436
rect 13817 14433 13829 14436
rect 13863 14433 13875 14467
rect 13817 14427 13875 14433
rect 13265 14399 13323 14405
rect 13265 14365 13277 14399
rect 13311 14365 13323 14399
rect 13265 14359 13323 14365
rect 13357 14399 13415 14405
rect 13357 14365 13369 14399
rect 13403 14365 13415 14399
rect 13357 14359 13415 14365
rect 13538 14356 13544 14408
rect 13596 14356 13602 14408
rect 13630 14356 13636 14408
rect 13688 14356 13694 14408
rect 14292 14405 14320 14504
rect 14691 14501 14703 14504
rect 14737 14532 14749 14535
rect 15488 14532 15516 14572
rect 15565 14569 15577 14603
rect 15611 14600 15623 14603
rect 15654 14600 15660 14612
rect 15611 14572 15660 14600
rect 15611 14569 15623 14572
rect 15565 14563 15623 14569
rect 15654 14560 15660 14572
rect 15712 14560 15718 14612
rect 17126 14600 17132 14612
rect 16960 14572 17132 14600
rect 16960 14541 16988 14572
rect 17126 14560 17132 14572
rect 17184 14560 17190 14612
rect 24854 14560 24860 14612
rect 24912 14600 24918 14612
rect 25406 14600 25412 14612
rect 24912 14572 25412 14600
rect 24912 14560 24918 14572
rect 25406 14560 25412 14572
rect 25464 14600 25470 14612
rect 27617 14603 27675 14609
rect 27617 14600 27629 14603
rect 25464 14572 27629 14600
rect 25464 14560 25470 14572
rect 27617 14569 27629 14572
rect 27663 14569 27675 14603
rect 27617 14563 27675 14569
rect 15749 14535 15807 14541
rect 15749 14532 15761 14535
rect 14737 14504 15332 14532
rect 15488 14504 15761 14532
rect 14737 14501 14749 14504
rect 14691 14495 14749 14501
rect 15197 14467 15255 14473
rect 15197 14464 15209 14467
rect 14476 14436 15209 14464
rect 14476 14405 14504 14436
rect 14844 14408 14872 14436
rect 15197 14433 15209 14436
rect 15243 14433 15255 14467
rect 15197 14427 15255 14433
rect 15304 14408 15332 14504
rect 15749 14501 15761 14504
rect 15795 14501 15807 14535
rect 15749 14495 15807 14501
rect 16945 14535 17003 14541
rect 16945 14501 16957 14535
rect 16991 14501 17003 14535
rect 16945 14495 17003 14501
rect 23750 14492 23756 14544
rect 23808 14532 23814 14544
rect 24762 14532 24768 14544
rect 23808 14504 24768 14532
rect 23808 14492 23814 14504
rect 24762 14492 24768 14504
rect 24820 14532 24826 14544
rect 25317 14535 25375 14541
rect 25317 14532 25329 14535
rect 24820 14504 25329 14532
rect 24820 14492 24826 14504
rect 25317 14501 25329 14504
rect 25363 14501 25375 14535
rect 25317 14495 25375 14501
rect 17034 14424 17040 14476
rect 17092 14424 17098 14476
rect 17129 14467 17187 14473
rect 17129 14433 17141 14467
rect 17175 14464 17187 14467
rect 17218 14464 17224 14476
rect 17175 14436 17224 14464
rect 17175 14433 17187 14436
rect 17129 14427 17187 14433
rect 17218 14424 17224 14436
rect 17276 14424 17282 14476
rect 19150 14424 19156 14476
rect 19208 14464 19214 14476
rect 20714 14464 20720 14476
rect 19208 14436 20720 14464
rect 19208 14424 19214 14436
rect 20714 14424 20720 14436
rect 20772 14424 20778 14476
rect 22370 14424 22376 14476
rect 22428 14464 22434 14476
rect 24489 14467 24547 14473
rect 24489 14464 24501 14467
rect 22428 14436 24501 14464
rect 22428 14424 22434 14436
rect 24489 14433 24501 14436
rect 24535 14464 24547 14467
rect 25130 14464 25136 14476
rect 24535 14436 25136 14464
rect 24535 14433 24547 14436
rect 24489 14427 24547 14433
rect 25130 14424 25136 14436
rect 25188 14424 25194 14476
rect 13725 14399 13783 14405
rect 13725 14365 13737 14399
rect 13771 14365 13783 14399
rect 13725 14359 13783 14365
rect 14277 14399 14335 14405
rect 14277 14365 14289 14399
rect 14323 14365 14335 14399
rect 14277 14359 14335 14365
rect 14461 14399 14519 14405
rect 14461 14365 14473 14399
rect 14507 14365 14519 14399
rect 14461 14359 14519 14365
rect 14553 14399 14611 14405
rect 14553 14365 14565 14399
rect 14599 14396 14611 14399
rect 14599 14368 14780 14396
rect 14599 14365 14611 14368
rect 14553 14359 14611 14365
rect 11517 14331 11575 14337
rect 11517 14297 11529 14331
rect 11563 14297 11575 14331
rect 12894 14328 12900 14340
rect 12742 14300 12900 14328
rect 11517 14291 11575 14297
rect 2314 14220 2320 14272
rect 2372 14260 2378 14272
rect 3694 14260 3700 14272
rect 2372 14232 3700 14260
rect 2372 14220 2378 14232
rect 3694 14220 3700 14232
rect 3752 14220 3758 14272
rect 11532 14260 11560 14291
rect 12894 14288 12900 14300
rect 12952 14288 12958 14340
rect 13740 14328 13768 14359
rect 13004 14300 13768 14328
rect 13004 14272 13032 14300
rect 12250 14260 12256 14272
rect 11532 14232 12256 14260
rect 12250 14220 12256 14232
rect 12308 14220 12314 14272
rect 12986 14220 12992 14272
rect 13044 14220 13050 14272
rect 14369 14263 14427 14269
rect 14369 14229 14381 14263
rect 14415 14260 14427 14263
rect 14642 14260 14648 14272
rect 14415 14232 14648 14260
rect 14415 14229 14427 14232
rect 14369 14223 14427 14229
rect 14642 14220 14648 14232
rect 14700 14220 14706 14272
rect 14752 14260 14780 14368
rect 14826 14356 14832 14408
rect 14884 14356 14890 14408
rect 15010 14356 15016 14408
rect 15068 14356 15074 14408
rect 15105 14399 15163 14405
rect 15105 14365 15117 14399
rect 15151 14396 15163 14399
rect 15286 14396 15292 14408
rect 15151 14368 15292 14396
rect 15151 14365 15163 14368
rect 15105 14359 15163 14365
rect 15286 14356 15292 14368
rect 15344 14356 15350 14408
rect 15381 14399 15439 14405
rect 15381 14365 15393 14399
rect 15427 14396 15439 14399
rect 15654 14396 15660 14408
rect 15427 14368 15660 14396
rect 15427 14365 15439 14368
rect 15381 14359 15439 14365
rect 15654 14356 15660 14368
rect 15712 14356 15718 14408
rect 15948 14368 16528 14396
rect 14921 14331 14979 14337
rect 14921 14297 14933 14331
rect 14967 14328 14979 14331
rect 15948 14328 15976 14368
rect 14967 14300 15976 14328
rect 16025 14331 16083 14337
rect 14967 14297 14979 14300
rect 14921 14291 14979 14297
rect 16025 14297 16037 14331
rect 16071 14297 16083 14331
rect 16500 14328 16528 14368
rect 16666 14356 16672 14408
rect 16724 14356 16730 14408
rect 16758 14356 16764 14408
rect 16816 14356 16822 14408
rect 16945 14399 17003 14405
rect 16945 14365 16957 14399
rect 16991 14396 17003 14399
rect 17862 14396 17868 14408
rect 16991 14368 17868 14396
rect 16991 14365 17003 14368
rect 16945 14359 17003 14365
rect 17862 14356 17868 14368
rect 17920 14356 17926 14408
rect 18414 14356 18420 14408
rect 18472 14396 18478 14408
rect 19058 14396 19064 14408
rect 18472 14368 19064 14396
rect 18472 14356 18478 14368
rect 19058 14356 19064 14368
rect 19116 14396 19122 14408
rect 20349 14399 20407 14405
rect 20349 14396 20361 14399
rect 19116 14368 20361 14396
rect 19116 14356 19122 14368
rect 20349 14365 20361 14368
rect 20395 14396 20407 14399
rect 20395 14368 22094 14396
rect 20395 14365 20407 14368
rect 20349 14359 20407 14365
rect 18230 14328 18236 14340
rect 16500 14300 18236 14328
rect 16025 14291 16083 14297
rect 15654 14260 15660 14272
rect 14752 14232 15660 14260
rect 15654 14220 15660 14232
rect 15712 14220 15718 14272
rect 16040 14260 16068 14291
rect 18230 14288 18236 14300
rect 18288 14288 18294 14340
rect 18432 14260 18460 14356
rect 19702 14288 19708 14340
rect 19760 14328 19766 14340
rect 20622 14328 20628 14340
rect 19760 14300 20628 14328
rect 19760 14288 19766 14300
rect 20622 14288 20628 14300
rect 20680 14288 20686 14340
rect 22066 14328 22094 14368
rect 24578 14356 24584 14408
rect 24636 14356 24642 14408
rect 27798 14356 27804 14408
rect 27856 14356 27862 14408
rect 22066 14300 22968 14328
rect 16040 14232 18460 14260
rect 20257 14263 20315 14269
rect 20257 14229 20269 14263
rect 20303 14260 20315 14263
rect 20438 14260 20444 14272
rect 20303 14232 20444 14260
rect 20303 14229 20315 14232
rect 20257 14223 20315 14229
rect 20438 14220 20444 14232
rect 20496 14220 20502 14272
rect 20530 14220 20536 14272
rect 20588 14260 20594 14272
rect 22830 14260 22836 14272
rect 20588 14232 22836 14260
rect 20588 14220 20594 14232
rect 22830 14220 22836 14232
rect 22888 14220 22894 14272
rect 22940 14260 22968 14300
rect 23290 14288 23296 14340
rect 23348 14288 23354 14340
rect 24118 14288 24124 14340
rect 24176 14328 24182 14340
rect 25133 14331 25191 14337
rect 25133 14328 25145 14331
rect 24176 14300 25145 14328
rect 24176 14288 24182 14300
rect 25133 14297 25145 14300
rect 25179 14297 25191 14331
rect 25133 14291 25191 14297
rect 23569 14263 23627 14269
rect 23569 14260 23581 14263
rect 22940 14232 23581 14260
rect 23569 14229 23581 14232
rect 23615 14260 23627 14263
rect 23842 14260 23848 14272
rect 23615 14232 23848 14260
rect 23615 14229 23627 14232
rect 23569 14223 23627 14229
rect 23842 14220 23848 14232
rect 23900 14220 23906 14272
rect 24946 14220 24952 14272
rect 25004 14220 25010 14272
rect 1104 14170 28152 14192
rect 1104 14118 4874 14170
rect 4926 14118 4938 14170
rect 4990 14118 5002 14170
rect 5054 14118 5066 14170
rect 5118 14118 5130 14170
rect 5182 14118 28152 14170
rect 1104 14096 28152 14118
rect 2774 14016 2780 14068
rect 2832 14056 2838 14068
rect 2832 14028 3556 14056
rect 2832 14016 2838 14028
rect 1673 13991 1731 13997
rect 1673 13957 1685 13991
rect 1719 13988 1731 13991
rect 1719 13960 2728 13988
rect 1719 13957 1731 13960
rect 1673 13951 1731 13957
rect 2700 13932 2728 13960
rect 3234 13948 3240 14000
rect 3292 13948 3298 14000
rect 1394 13880 1400 13932
rect 1452 13880 1458 13932
rect 2225 13923 2283 13929
rect 2225 13889 2237 13923
rect 2271 13889 2283 13923
rect 2225 13883 2283 13889
rect 2240 13796 2268 13883
rect 2682 13880 2688 13932
rect 2740 13920 2746 13932
rect 3053 13923 3111 13929
rect 3053 13920 3065 13923
rect 2740 13892 3065 13920
rect 2740 13880 2746 13892
rect 3053 13889 3065 13892
rect 3099 13889 3111 13923
rect 3053 13883 3111 13889
rect 3142 13880 3148 13932
rect 3200 13880 3206 13932
rect 3252 13920 3280 13948
rect 3421 13923 3479 13929
rect 3421 13920 3433 13923
rect 3252 13892 3433 13920
rect 3421 13889 3433 13892
rect 3467 13889 3479 13923
rect 3528 13920 3556 14028
rect 3602 14016 3608 14068
rect 3660 14016 3666 14068
rect 16482 14056 16488 14068
rect 11532 14028 16488 14056
rect 3605 13923 3663 13929
rect 3605 13920 3617 13923
rect 3528 13892 3617 13920
rect 3421 13883 3479 13889
rect 3605 13889 3617 13892
rect 3651 13889 3663 13923
rect 3605 13883 3663 13889
rect 3694 13880 3700 13932
rect 3752 13880 3758 13932
rect 3881 13923 3939 13929
rect 3881 13889 3893 13923
rect 3927 13889 3939 13923
rect 3881 13883 3939 13889
rect 2314 13812 2320 13864
rect 2372 13812 2378 13864
rect 2593 13855 2651 13861
rect 2593 13821 2605 13855
rect 2639 13852 2651 13855
rect 2958 13852 2964 13864
rect 2639 13824 2964 13852
rect 2639 13821 2651 13824
rect 2593 13815 2651 13821
rect 2958 13812 2964 13824
rect 3016 13812 3022 13864
rect 3237 13855 3295 13861
rect 3237 13821 3249 13855
rect 3283 13852 3295 13855
rect 3789 13855 3847 13861
rect 3789 13852 3801 13855
rect 3283 13824 3801 13852
rect 3283 13821 3295 13824
rect 3237 13815 3295 13821
rect 3789 13821 3801 13824
rect 3835 13821 3847 13855
rect 3789 13815 3847 13821
rect 2222 13744 2228 13796
rect 2280 13784 2286 13796
rect 3896 13784 3924 13883
rect 4154 13880 4160 13932
rect 4212 13880 4218 13932
rect 4246 13880 4252 13932
rect 4304 13920 4310 13932
rect 4341 13923 4399 13929
rect 4341 13920 4353 13923
rect 4304 13892 4353 13920
rect 4304 13880 4310 13892
rect 4341 13889 4353 13892
rect 4387 13920 4399 13923
rect 4798 13920 4804 13932
rect 4387 13892 4804 13920
rect 4387 13889 4399 13892
rect 4341 13883 4399 13889
rect 4798 13880 4804 13892
rect 4856 13880 4862 13932
rect 5813 13923 5871 13929
rect 5813 13889 5825 13923
rect 5859 13920 5871 13923
rect 6730 13920 6736 13932
rect 5859 13892 6736 13920
rect 5859 13889 5871 13892
rect 5813 13883 5871 13889
rect 6730 13880 6736 13892
rect 6788 13880 6794 13932
rect 6917 13923 6975 13929
rect 6917 13889 6929 13923
rect 6963 13889 6975 13923
rect 6917 13883 6975 13889
rect 5902 13812 5908 13864
rect 5960 13812 5966 13864
rect 6932 13796 6960 13883
rect 7006 13880 7012 13932
rect 7064 13920 7070 13932
rect 7193 13923 7251 13929
rect 7193 13920 7205 13923
rect 7064 13892 7205 13920
rect 7064 13880 7070 13892
rect 7193 13889 7205 13892
rect 7239 13889 7251 13923
rect 7193 13883 7251 13889
rect 7558 13880 7564 13932
rect 7616 13880 7622 13932
rect 8294 13880 8300 13932
rect 8352 13920 8358 13932
rect 9401 13923 9459 13929
rect 9401 13920 9413 13923
rect 8352 13892 9413 13920
rect 8352 13880 8358 13892
rect 9401 13889 9413 13892
rect 9447 13889 9459 13923
rect 9401 13883 9459 13889
rect 9582 13880 9588 13932
rect 9640 13880 9646 13932
rect 9674 13880 9680 13932
rect 9732 13880 9738 13932
rect 11238 13880 11244 13932
rect 11296 13920 11302 13932
rect 11532 13929 11560 14028
rect 11793 13991 11851 13997
rect 11793 13957 11805 13991
rect 11839 13988 11851 13991
rect 11882 13988 11888 14000
rect 11839 13960 11888 13988
rect 11839 13957 11851 13960
rect 11793 13951 11851 13957
rect 11882 13948 11888 13960
rect 11940 13948 11946 14000
rect 13446 13948 13452 14000
rect 13504 13948 13510 14000
rect 11517 13923 11575 13929
rect 11517 13920 11529 13923
rect 11296 13892 11529 13920
rect 11296 13880 11302 13892
rect 11517 13889 11529 13892
rect 11563 13889 11575 13923
rect 11517 13883 11575 13889
rect 12894 13880 12900 13932
rect 12952 13880 12958 13932
rect 13078 13880 13084 13932
rect 13136 13920 13142 13932
rect 13725 13923 13783 13929
rect 13725 13920 13737 13923
rect 13136 13892 13737 13920
rect 13136 13880 13142 13892
rect 13725 13889 13737 13892
rect 13771 13889 13783 13923
rect 13725 13883 13783 13889
rect 14090 13880 14096 13932
rect 14148 13920 14154 13932
rect 14384 13929 14412 14028
rect 16482 14016 16488 14028
rect 16540 14016 16546 14068
rect 17126 14016 17132 14068
rect 17184 14056 17190 14068
rect 17405 14059 17463 14065
rect 17405 14056 17417 14059
rect 17184 14028 17417 14056
rect 17184 14016 17190 14028
rect 17405 14025 17417 14028
rect 17451 14025 17463 14059
rect 18598 14056 18604 14068
rect 17405 14019 17463 14025
rect 18340 14028 18604 14056
rect 14642 13948 14648 14000
rect 14700 13948 14706 14000
rect 16574 13988 16580 14000
rect 15870 13974 16580 13988
rect 15856 13960 16580 13974
rect 14185 13923 14243 13929
rect 14185 13920 14197 13923
rect 14148 13892 14197 13920
rect 14148 13880 14154 13892
rect 14185 13889 14197 13892
rect 14231 13889 14243 13923
rect 14185 13883 14243 13889
rect 14369 13923 14427 13929
rect 14369 13889 14381 13923
rect 14415 13889 14427 13923
rect 14369 13883 14427 13889
rect 8662 13812 8668 13864
rect 8720 13812 8726 13864
rect 12912 13852 12940 13880
rect 15856 13852 15884 13960
rect 16574 13948 16580 13960
rect 16632 13948 16638 14000
rect 17037 13991 17095 13997
rect 17037 13988 17049 13991
rect 16684 13960 17049 13988
rect 15930 13880 15936 13932
rect 15988 13920 15994 13932
rect 16684 13920 16712 13960
rect 17037 13957 17049 13960
rect 17083 13957 17095 13991
rect 17037 13951 17095 13957
rect 18049 13991 18107 13997
rect 18049 13957 18061 13991
rect 18095 13988 18107 13991
rect 18230 13988 18236 14000
rect 18095 13960 18236 13988
rect 18095 13957 18107 13960
rect 18049 13951 18107 13957
rect 18230 13948 18236 13960
rect 18288 13948 18294 14000
rect 15988 13892 16712 13920
rect 15988 13880 15994 13892
rect 16850 13880 16856 13932
rect 16908 13880 16914 13932
rect 17129 13923 17187 13929
rect 17129 13889 17141 13923
rect 17175 13889 17187 13923
rect 17129 13883 17187 13889
rect 17221 13923 17279 13929
rect 17221 13889 17233 13923
rect 17267 13920 17279 13923
rect 18340 13920 18368 14028
rect 18598 14016 18604 14028
rect 18656 14016 18662 14068
rect 19245 14059 19303 14065
rect 19245 14025 19257 14059
rect 19291 14056 19303 14059
rect 20530 14056 20536 14068
rect 19291 14028 20536 14056
rect 19291 14025 19303 14028
rect 19245 14019 19303 14025
rect 20530 14016 20536 14028
rect 20588 14016 20594 14068
rect 20714 14016 20720 14068
rect 20772 14056 20778 14068
rect 21542 14056 21548 14068
rect 20772 14028 21548 14056
rect 20772 14016 20778 14028
rect 21542 14016 21548 14028
rect 21600 14056 21606 14068
rect 23382 14056 23388 14068
rect 21600 14028 23388 14056
rect 21600 14016 21606 14028
rect 18414 13948 18420 14000
rect 18472 13948 18478 14000
rect 18874 13948 18880 14000
rect 18932 13988 18938 14000
rect 18932 13960 19104 13988
rect 18932 13948 18938 13960
rect 17267 13892 18368 13920
rect 17267 13889 17279 13892
rect 17221 13883 17279 13889
rect 12912 13824 15884 13852
rect 17144 13852 17172 13883
rect 17770 13852 17776 13864
rect 17144 13824 17776 13852
rect 17770 13812 17776 13824
rect 17828 13812 17834 13864
rect 17954 13812 17960 13864
rect 18012 13852 18018 13864
rect 18432 13861 18460 13948
rect 18601 13923 18659 13929
rect 18601 13889 18613 13923
rect 18647 13889 18659 13923
rect 18601 13883 18659 13889
rect 18693 13926 18751 13929
rect 18782 13926 18788 13932
rect 18693 13923 18788 13926
rect 18693 13889 18705 13923
rect 18739 13898 18788 13923
rect 18739 13889 18751 13898
rect 18693 13883 18751 13889
rect 18233 13855 18291 13861
rect 18012 13824 18184 13852
rect 18012 13812 18018 13824
rect 2280 13756 3924 13784
rect 6181 13787 6239 13793
rect 2280 13744 2286 13756
rect 6181 13753 6193 13787
rect 6227 13784 6239 13787
rect 6914 13784 6920 13796
rect 6227 13756 6920 13784
rect 6227 13753 6239 13756
rect 6181 13747 6239 13753
rect 6914 13744 6920 13756
rect 6972 13744 6978 13796
rect 7469 13787 7527 13793
rect 7469 13753 7481 13787
rect 7515 13784 7527 13787
rect 8570 13784 8576 13796
rect 7515 13756 8576 13784
rect 7515 13753 7527 13756
rect 7469 13747 7527 13753
rect 8570 13744 8576 13756
rect 8628 13784 8634 13796
rect 8941 13787 8999 13793
rect 8941 13784 8953 13787
rect 8628 13756 8953 13784
rect 8628 13744 8634 13756
rect 8941 13753 8953 13756
rect 8987 13753 8999 13787
rect 8941 13747 8999 13753
rect 13722 13744 13728 13796
rect 13780 13784 13786 13796
rect 18156 13793 18184 13824
rect 18233 13821 18245 13855
rect 18279 13821 18291 13855
rect 18233 13815 18291 13821
rect 18325 13855 18383 13861
rect 18325 13821 18337 13855
rect 18371 13821 18383 13855
rect 18325 13815 18383 13821
rect 18417 13855 18475 13861
rect 18417 13821 18429 13855
rect 18463 13821 18475 13855
rect 18616 13852 18644 13883
rect 18782 13880 18788 13898
rect 18840 13880 18846 13932
rect 18966 13880 18972 13932
rect 19024 13880 19030 13932
rect 19076 13929 19104 13960
rect 19150 13948 19156 14000
rect 19208 13988 19214 14000
rect 19981 13991 20039 13997
rect 19208 13960 19932 13988
rect 19208 13948 19214 13960
rect 19061 13923 19119 13929
rect 19061 13889 19073 13923
rect 19107 13889 19119 13923
rect 19061 13883 19119 13889
rect 19521 13923 19579 13929
rect 19521 13889 19533 13923
rect 19567 13920 19579 13923
rect 19702 13920 19708 13932
rect 19567 13892 19708 13920
rect 19567 13889 19579 13892
rect 19521 13883 19579 13889
rect 19702 13880 19708 13892
rect 19760 13880 19766 13932
rect 19797 13923 19855 13929
rect 19797 13889 19809 13923
rect 19843 13889 19855 13923
rect 19904 13920 19932 13960
rect 19981 13957 19993 13991
rect 20027 13988 20039 13991
rect 21085 13991 21143 13997
rect 21085 13988 21097 13991
rect 20027 13960 21097 13988
rect 20027 13957 20039 13960
rect 19981 13951 20039 13957
rect 20364 13929 20392 13960
rect 21085 13957 21097 13960
rect 21131 13957 21143 13991
rect 21358 13988 21364 14000
rect 21085 13951 21143 13957
rect 21192 13960 21364 13988
rect 20073 13923 20131 13929
rect 20073 13920 20085 13923
rect 19904 13892 20085 13920
rect 19797 13883 19855 13889
rect 20073 13889 20085 13892
rect 20119 13889 20131 13923
rect 20073 13883 20131 13889
rect 20338 13923 20396 13929
rect 20338 13889 20350 13923
rect 20384 13889 20396 13923
rect 20338 13883 20396 13889
rect 20717 13923 20775 13929
rect 20717 13889 20729 13923
rect 20763 13889 20775 13923
rect 20717 13883 20775 13889
rect 18874 13852 18880 13864
rect 18616 13824 18880 13852
rect 18417 13815 18475 13821
rect 14001 13787 14059 13793
rect 14001 13784 14013 13787
rect 13780 13756 14013 13784
rect 13780 13744 13786 13756
rect 14001 13753 14013 13756
rect 14047 13753 14059 13787
rect 14001 13747 14059 13753
rect 18141 13787 18199 13793
rect 18141 13753 18153 13787
rect 18187 13753 18199 13787
rect 18141 13747 18199 13753
rect 4341 13719 4399 13725
rect 4341 13685 4353 13719
rect 4387 13716 4399 13719
rect 4614 13716 4620 13728
rect 4387 13688 4620 13716
rect 4387 13685 4399 13688
rect 4341 13679 4399 13685
rect 4614 13676 4620 13688
rect 4672 13676 4678 13728
rect 9122 13676 9128 13728
rect 9180 13676 9186 13728
rect 9214 13676 9220 13728
rect 9272 13676 9278 13728
rect 12802 13676 12808 13728
rect 12860 13716 12866 13728
rect 13265 13719 13323 13725
rect 13265 13716 13277 13719
rect 12860 13688 13277 13716
rect 12860 13676 12866 13688
rect 13265 13685 13277 13688
rect 13311 13685 13323 13719
rect 13265 13679 13323 13685
rect 13814 13676 13820 13728
rect 13872 13676 13878 13728
rect 13909 13719 13967 13725
rect 13909 13685 13921 13719
rect 13955 13716 13967 13719
rect 14734 13716 14740 13728
rect 13955 13688 14740 13716
rect 13955 13685 13967 13688
rect 13909 13679 13967 13685
rect 14734 13676 14740 13688
rect 14792 13676 14798 13728
rect 15378 13676 15384 13728
rect 15436 13716 15442 13728
rect 16117 13719 16175 13725
rect 16117 13716 16129 13719
rect 15436 13688 16129 13716
rect 15436 13676 15442 13688
rect 16117 13685 16129 13688
rect 16163 13685 16175 13719
rect 16117 13679 16175 13685
rect 18046 13676 18052 13728
rect 18104 13716 18110 13728
rect 18248 13716 18276 13815
rect 18340 13784 18368 13815
rect 18874 13812 18880 13824
rect 18932 13852 18938 13864
rect 19429 13855 19487 13861
rect 19429 13852 19441 13855
rect 18932 13824 19441 13852
rect 18932 13812 18938 13824
rect 19429 13821 19441 13824
rect 19475 13821 19487 13855
rect 19812 13852 19840 13883
rect 20438 13852 20444 13864
rect 19812 13824 20444 13852
rect 19429 13815 19487 13821
rect 20438 13812 20444 13824
rect 20496 13812 20502 13864
rect 20530 13812 20536 13864
rect 20588 13812 20594 13864
rect 20622 13812 20628 13864
rect 20680 13812 20686 13864
rect 20732 13852 20760 13883
rect 20898 13880 20904 13932
rect 20956 13880 20962 13932
rect 21192 13929 21220 13960
rect 21358 13948 21364 13960
rect 21416 13948 21422 14000
rect 21453 13991 21511 13997
rect 21453 13957 21465 13991
rect 21499 13988 21511 13991
rect 22370 13988 22376 14000
rect 21499 13960 22376 13988
rect 21499 13957 21511 13960
rect 21453 13951 21511 13957
rect 22370 13948 22376 13960
rect 22428 13948 22434 14000
rect 21177 13923 21235 13929
rect 21177 13889 21189 13923
rect 21223 13889 21235 13923
rect 21177 13883 21235 13889
rect 21634 13880 21640 13932
rect 21692 13880 21698 13932
rect 22189 13923 22247 13929
rect 22189 13889 22201 13923
rect 22235 13889 22247 13923
rect 22189 13883 22247 13889
rect 21269 13855 21327 13861
rect 21269 13852 21281 13855
rect 20732 13824 21281 13852
rect 21269 13821 21281 13824
rect 21315 13821 21327 13855
rect 22204 13852 22232 13883
rect 22278 13880 22284 13932
rect 22336 13880 22342 13932
rect 22462 13880 22468 13932
rect 22520 13880 22526 13932
rect 22554 13880 22560 13932
rect 22612 13880 22618 13932
rect 22664 13920 22692 14028
rect 23382 14016 23388 14028
rect 23440 14016 23446 14068
rect 24578 14016 24584 14068
rect 24636 14056 24642 14068
rect 25685 14059 25743 14065
rect 25685 14056 25697 14059
rect 24636 14028 25697 14056
rect 24636 14016 24642 14028
rect 25685 14025 25697 14028
rect 25731 14025 25743 14059
rect 25685 14019 25743 14025
rect 22741 13991 22799 13997
rect 22741 13957 22753 13991
rect 22787 13988 22799 13991
rect 22787 13960 23428 13988
rect 22787 13957 22799 13960
rect 22741 13951 22799 13957
rect 22833 13923 22891 13929
rect 22833 13920 22845 13923
rect 22664 13892 22845 13920
rect 22833 13889 22845 13892
rect 22879 13889 22891 13923
rect 22833 13883 22891 13889
rect 23014 13880 23020 13932
rect 23072 13880 23078 13932
rect 23400 13929 23428 13960
rect 25222 13948 25228 14000
rect 25280 13948 25286 14000
rect 23385 13923 23443 13929
rect 23385 13889 23397 13923
rect 23431 13889 23443 13923
rect 23385 13883 23443 13889
rect 23474 13880 23480 13932
rect 23532 13920 23538 13932
rect 23937 13923 23995 13929
rect 23937 13920 23949 13923
rect 23532 13892 23949 13920
rect 23532 13880 23538 13892
rect 23937 13889 23949 13892
rect 23983 13889 23995 13923
rect 23937 13883 23995 13889
rect 23032 13852 23060 13880
rect 22204 13824 23060 13852
rect 21269 13815 21327 13821
rect 23566 13812 23572 13864
rect 23624 13812 23630 13864
rect 23842 13812 23848 13864
rect 23900 13812 23906 13864
rect 24213 13855 24271 13861
rect 24213 13852 24225 13855
rect 24044 13824 24225 13852
rect 18340 13756 18460 13784
rect 18104 13688 18276 13716
rect 18432 13716 18460 13756
rect 18598 13744 18604 13796
rect 18656 13784 18662 13796
rect 18785 13787 18843 13793
rect 18785 13784 18797 13787
rect 18656 13756 18797 13784
rect 18656 13744 18662 13756
rect 18785 13753 18797 13756
rect 18831 13784 18843 13787
rect 18831 13756 19334 13784
rect 18831 13753 18843 13756
rect 18785 13747 18843 13753
rect 18966 13716 18972 13728
rect 18432 13688 18972 13716
rect 18104 13676 18110 13688
rect 18966 13676 18972 13688
rect 19024 13676 19030 13728
rect 19306 13716 19334 13756
rect 20254 13744 20260 13796
rect 20312 13784 20318 13796
rect 22554 13784 22560 13796
rect 20312 13756 22560 13784
rect 20312 13744 20318 13756
rect 22554 13744 22560 13756
rect 22612 13744 22618 13796
rect 22922 13744 22928 13796
rect 22980 13784 22986 13796
rect 23753 13787 23811 13793
rect 23753 13784 23765 13787
rect 22980 13756 23765 13784
rect 22980 13744 22986 13756
rect 23753 13753 23765 13756
rect 23799 13784 23811 13787
rect 24044 13784 24072 13824
rect 24213 13821 24225 13824
rect 24259 13821 24271 13855
rect 24213 13815 24271 13821
rect 23799 13756 24072 13784
rect 23799 13753 23811 13756
rect 23753 13747 23811 13753
rect 19518 13716 19524 13728
rect 19306 13688 19524 13716
rect 19518 13676 19524 13688
rect 19576 13676 19582 13728
rect 19610 13676 19616 13728
rect 19668 13676 19674 13728
rect 19978 13676 19984 13728
rect 20036 13716 20042 13728
rect 20165 13719 20223 13725
rect 20165 13716 20177 13719
rect 20036 13688 20177 13716
rect 20036 13676 20042 13688
rect 20165 13685 20177 13688
rect 20211 13685 20223 13719
rect 20165 13679 20223 13685
rect 20346 13676 20352 13728
rect 20404 13716 20410 13728
rect 23382 13716 23388 13728
rect 20404 13688 23388 13716
rect 20404 13676 20410 13688
rect 23382 13676 23388 13688
rect 23440 13676 23446 13728
rect 1104 13626 28152 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 28152 13626
rect 1104 13552 28152 13574
rect 4908 13484 8248 13512
rect 4908 13444 4936 13484
rect 8220 13456 8248 13484
rect 8754 13472 8760 13524
rect 8812 13472 8818 13524
rect 10226 13472 10232 13524
rect 10284 13512 10290 13524
rect 10410 13512 10416 13524
rect 10284 13484 10416 13512
rect 10284 13472 10290 13484
rect 10410 13472 10416 13484
rect 10468 13472 10474 13524
rect 12989 13515 13047 13521
rect 12989 13481 13001 13515
rect 13035 13512 13047 13515
rect 13814 13512 13820 13524
rect 13035 13484 13820 13512
rect 13035 13481 13047 13484
rect 12989 13475 13047 13481
rect 13814 13472 13820 13484
rect 13872 13472 13878 13524
rect 14826 13472 14832 13524
rect 14884 13512 14890 13524
rect 14921 13515 14979 13521
rect 14921 13512 14933 13515
rect 14884 13484 14933 13512
rect 14884 13472 14890 13484
rect 14921 13481 14933 13484
rect 14967 13481 14979 13515
rect 14921 13475 14979 13481
rect 15286 13472 15292 13524
rect 15344 13512 15350 13524
rect 15473 13515 15531 13521
rect 15473 13512 15485 13515
rect 15344 13484 15485 13512
rect 15344 13472 15350 13484
rect 15473 13481 15485 13484
rect 15519 13481 15531 13515
rect 15473 13475 15531 13481
rect 15562 13472 15568 13524
rect 15620 13512 15626 13524
rect 15838 13512 15844 13524
rect 15620 13484 15844 13512
rect 15620 13472 15626 13484
rect 15838 13472 15844 13484
rect 15896 13472 15902 13524
rect 18509 13515 18567 13521
rect 18509 13481 18521 13515
rect 18555 13512 18567 13515
rect 18966 13512 18972 13524
rect 18555 13484 18972 13512
rect 18555 13481 18567 13484
rect 18509 13475 18567 13481
rect 18966 13472 18972 13484
rect 19024 13512 19030 13524
rect 19610 13512 19616 13524
rect 19024 13484 19616 13512
rect 19024 13472 19030 13484
rect 19610 13472 19616 13484
rect 19668 13472 19674 13524
rect 19702 13472 19708 13524
rect 19760 13512 19766 13524
rect 20346 13512 20352 13524
rect 19760 13484 20352 13512
rect 19760 13472 19766 13484
rect 20346 13472 20352 13484
rect 20404 13472 20410 13524
rect 21358 13472 21364 13524
rect 21416 13512 21422 13524
rect 21453 13515 21511 13521
rect 21453 13512 21465 13515
rect 21416 13484 21465 13512
rect 21416 13472 21422 13484
rect 21453 13481 21465 13484
rect 21499 13481 21511 13515
rect 21453 13475 21511 13481
rect 21545 13515 21603 13521
rect 21545 13481 21557 13515
rect 21591 13512 21603 13515
rect 21634 13512 21640 13524
rect 21591 13484 21640 13512
rect 21591 13481 21603 13484
rect 21545 13475 21603 13481
rect 2746 13416 4936 13444
rect 6917 13447 6975 13453
rect 2746 13252 2774 13416
rect 2958 13336 2964 13388
rect 3016 13336 3022 13388
rect 2869 13311 2927 13317
rect 2869 13277 2881 13311
rect 2915 13277 2927 13311
rect 2869 13271 2927 13277
rect 2682 13200 2688 13252
rect 2740 13212 2774 13252
rect 2884 13240 2912 13271
rect 3142 13268 3148 13320
rect 3200 13308 3206 13320
rect 3528 13317 3556 13416
rect 6917 13413 6929 13447
rect 6963 13413 6975 13447
rect 6917 13407 6975 13413
rect 4706 13336 4712 13388
rect 4764 13336 4770 13388
rect 6932 13376 6960 13407
rect 8202 13404 8208 13456
rect 8260 13444 8266 13456
rect 13173 13447 13231 13453
rect 8260 13416 9352 13444
rect 8260 13404 8266 13416
rect 8662 13376 8668 13388
rect 6932 13348 8668 13376
rect 3329 13311 3387 13317
rect 3329 13308 3341 13311
rect 3200 13280 3341 13308
rect 3200 13268 3206 13280
rect 3329 13277 3341 13280
rect 3375 13277 3387 13311
rect 3329 13271 3387 13277
rect 3513 13311 3571 13317
rect 3513 13277 3525 13311
rect 3559 13277 3571 13311
rect 3513 13271 3571 13277
rect 4614 13268 4620 13320
rect 4672 13268 4678 13320
rect 6914 13268 6920 13320
rect 6972 13268 6978 13320
rect 7006 13268 7012 13320
rect 7064 13308 7070 13320
rect 7193 13311 7251 13317
rect 7193 13308 7205 13311
rect 7064 13280 7205 13308
rect 7064 13268 7070 13280
rect 7193 13277 7205 13280
rect 7239 13277 7251 13311
rect 7193 13271 7251 13277
rect 8202 13268 8208 13320
rect 8260 13268 8266 13320
rect 8312 13317 8340 13348
rect 8662 13336 8668 13348
rect 8720 13336 8726 13388
rect 9122 13336 9128 13388
rect 9180 13336 9186 13388
rect 8297 13311 8355 13317
rect 8297 13277 8309 13311
rect 8343 13277 8355 13311
rect 8297 13271 8355 13277
rect 8478 13268 8484 13320
rect 8536 13268 8542 13320
rect 8573 13311 8631 13317
rect 8573 13277 8585 13311
rect 8619 13277 8631 13311
rect 8573 13271 8631 13277
rect 3421 13243 3479 13249
rect 3421 13240 3433 13243
rect 2884 13212 3433 13240
rect 2740 13200 2746 13212
rect 3421 13209 3433 13212
rect 3467 13209 3479 13243
rect 3421 13203 3479 13209
rect 7098 13200 7104 13252
rect 7156 13240 7162 13252
rect 7558 13240 7564 13252
rect 7156 13212 7564 13240
rect 7156 13200 7162 13212
rect 7558 13200 7564 13212
rect 7616 13200 7622 13252
rect 8588 13240 8616 13271
rect 9214 13268 9220 13320
rect 9272 13268 9278 13320
rect 9324 13308 9352 13416
rect 13173 13413 13185 13447
rect 13219 13444 13231 13447
rect 17034 13444 17040 13456
rect 13219 13416 17040 13444
rect 13219 13413 13231 13416
rect 13173 13407 13231 13413
rect 17034 13404 17040 13416
rect 17092 13404 17098 13456
rect 18601 13447 18659 13453
rect 18601 13413 18613 13447
rect 18647 13413 18659 13447
rect 18601 13407 18659 13413
rect 12069 13379 12127 13385
rect 12069 13345 12081 13379
rect 12115 13376 12127 13379
rect 12250 13376 12256 13388
rect 12115 13348 12256 13376
rect 12115 13345 12127 13348
rect 12069 13339 12127 13345
rect 12250 13336 12256 13348
rect 12308 13376 12314 13388
rect 13906 13376 13912 13388
rect 12308 13348 13124 13376
rect 12308 13336 12314 13348
rect 10137 13311 10195 13317
rect 10137 13308 10149 13311
rect 9324 13280 10149 13308
rect 10137 13277 10149 13280
rect 10183 13308 10195 13311
rect 10226 13308 10232 13320
rect 10183 13280 10232 13308
rect 10183 13277 10195 13280
rect 10137 13271 10195 13277
rect 10226 13268 10232 13280
rect 10284 13268 10290 13320
rect 11977 13311 12035 13317
rect 11977 13277 11989 13311
rect 12023 13308 12035 13311
rect 12342 13308 12348 13320
rect 12023 13280 12348 13308
rect 12023 13277 12035 13280
rect 11977 13271 12035 13277
rect 12342 13268 12348 13280
rect 12400 13268 12406 13320
rect 12710 13268 12716 13320
rect 12768 13268 12774 13320
rect 12802 13268 12808 13320
rect 12860 13268 12866 13320
rect 12986 13268 12992 13320
rect 13044 13268 13050 13320
rect 13096 13317 13124 13348
rect 13188 13348 13912 13376
rect 13081 13311 13139 13317
rect 13081 13277 13093 13311
rect 13127 13277 13139 13311
rect 13081 13271 13139 13277
rect 9674 13240 9680 13252
rect 8588 13212 9680 13240
rect 9674 13200 9680 13212
rect 9732 13200 9738 13252
rect 11609 13243 11667 13249
rect 11609 13209 11621 13243
rect 11655 13209 11667 13243
rect 11609 13203 11667 13209
rect 3237 13175 3295 13181
rect 3237 13141 3249 13175
rect 3283 13172 3295 13175
rect 3786 13172 3792 13184
rect 3283 13144 3792 13172
rect 3283 13141 3295 13144
rect 3237 13135 3295 13141
rect 3786 13132 3792 13144
rect 3844 13132 3850 13184
rect 5258 13132 5264 13184
rect 5316 13132 5322 13184
rect 10042 13132 10048 13184
rect 10100 13132 10106 13184
rect 11624 13172 11652 13203
rect 11698 13200 11704 13252
rect 11756 13200 11762 13252
rect 13188 13240 13216 13348
rect 13906 13336 13912 13348
rect 13964 13336 13970 13388
rect 13998 13336 14004 13388
rect 14056 13376 14062 13388
rect 15304 13376 15516 13384
rect 14056 13356 15516 13376
rect 14056 13348 15332 13356
rect 14056 13336 14062 13348
rect 13265 13311 13323 13317
rect 13265 13277 13277 13311
rect 13311 13277 13323 13311
rect 13265 13271 13323 13277
rect 12406 13212 13216 13240
rect 12158 13172 12164 13184
rect 11624 13144 12164 13172
rect 12158 13132 12164 13144
rect 12216 13132 12222 13184
rect 12253 13175 12311 13181
rect 12253 13141 12265 13175
rect 12299 13172 12311 13175
rect 12406 13172 12434 13212
rect 12299 13144 12434 13172
rect 12299 13141 12311 13144
rect 12253 13135 12311 13141
rect 12526 13132 12532 13184
rect 12584 13172 12590 13184
rect 13280 13172 13308 13271
rect 13538 13268 13544 13320
rect 13596 13268 13602 13320
rect 14642 13268 14648 13320
rect 14700 13268 14706 13320
rect 14829 13311 14887 13317
rect 14829 13277 14841 13311
rect 14875 13308 14887 13311
rect 14918 13308 14924 13320
rect 14875 13280 14924 13308
rect 14875 13277 14887 13280
rect 14829 13271 14887 13277
rect 14918 13268 14924 13280
rect 14976 13268 14982 13320
rect 15102 13268 15108 13320
rect 15160 13268 15166 13320
rect 15286 13268 15292 13320
rect 15344 13268 15350 13320
rect 15381 13311 15439 13317
rect 15381 13277 15393 13311
rect 15427 13307 15439 13311
rect 15488 13307 15516 13356
rect 15838 13336 15844 13388
rect 15896 13336 15902 13388
rect 15930 13336 15936 13388
rect 15988 13336 15994 13388
rect 16669 13379 16727 13385
rect 16669 13376 16681 13379
rect 16040 13348 16681 13376
rect 15427 13279 15516 13307
rect 15427 13277 15439 13279
rect 15381 13271 15439 13277
rect 15654 13268 15660 13320
rect 15712 13268 15718 13320
rect 16040 13317 16068 13348
rect 16669 13345 16681 13348
rect 16715 13345 16727 13379
rect 16669 13339 16727 13345
rect 17954 13336 17960 13388
rect 18012 13376 18018 13388
rect 18616 13376 18644 13407
rect 18012 13348 18644 13376
rect 18693 13379 18751 13385
rect 18012 13336 18018 13348
rect 18693 13345 18705 13379
rect 18739 13376 18751 13379
rect 18874 13376 18880 13388
rect 18739 13348 18880 13376
rect 18739 13345 18751 13348
rect 18693 13339 18751 13345
rect 18874 13336 18880 13348
rect 18932 13336 18938 13388
rect 19978 13376 19984 13388
rect 19444 13348 19984 13376
rect 16025 13311 16083 13317
rect 16025 13277 16037 13311
rect 16071 13277 16083 13311
rect 16025 13271 16083 13277
rect 16209 13311 16267 13317
rect 16209 13277 16221 13311
rect 16255 13308 16267 13311
rect 16255 13280 16712 13308
rect 16255 13277 16267 13280
rect 16209 13271 16267 13277
rect 14737 13243 14795 13249
rect 14737 13209 14749 13243
rect 14783 13240 14795 13243
rect 16301 13243 16359 13249
rect 16301 13240 16313 13243
rect 14783 13212 15240 13240
rect 14783 13209 14795 13212
rect 14737 13203 14795 13209
rect 13354 13172 13360 13184
rect 12584 13144 13360 13172
rect 12584 13132 12590 13144
rect 13354 13132 13360 13144
rect 13412 13132 13418 13184
rect 13725 13175 13783 13181
rect 13725 13141 13737 13175
rect 13771 13172 13783 13175
rect 14090 13172 14096 13184
rect 13771 13144 14096 13172
rect 13771 13141 13783 13144
rect 13725 13135 13783 13141
rect 14090 13132 14096 13144
rect 14148 13132 14154 13184
rect 15212 13172 15240 13212
rect 15488 13212 16313 13240
rect 15488 13172 15516 13212
rect 16301 13209 16313 13212
rect 16347 13209 16359 13243
rect 16301 13203 16359 13209
rect 16390 13200 16396 13252
rect 16448 13240 16454 13252
rect 16485 13243 16543 13249
rect 16485 13240 16497 13243
rect 16448 13212 16497 13240
rect 16448 13200 16454 13212
rect 16485 13209 16497 13212
rect 16531 13209 16543 13243
rect 16684 13240 16712 13280
rect 18414 13268 18420 13320
rect 18472 13308 18478 13320
rect 19444 13317 19472 13348
rect 19978 13336 19984 13348
rect 20036 13336 20042 13388
rect 21174 13336 21180 13388
rect 21232 13376 21238 13388
rect 21468 13376 21496 13475
rect 21634 13472 21640 13484
rect 21692 13472 21698 13524
rect 21726 13472 21732 13524
rect 21784 13512 21790 13524
rect 22186 13512 22192 13524
rect 21784 13484 22192 13512
rect 21784 13472 21790 13484
rect 22186 13472 22192 13484
rect 22244 13472 22250 13524
rect 22373 13515 22431 13521
rect 22373 13481 22385 13515
rect 22419 13512 22431 13515
rect 23290 13512 23296 13524
rect 22419 13484 23296 13512
rect 22419 13481 22431 13484
rect 22373 13475 22431 13481
rect 23290 13472 23296 13484
rect 23348 13472 23354 13524
rect 23566 13472 23572 13524
rect 23624 13512 23630 13524
rect 24397 13515 24455 13521
rect 24397 13512 24409 13515
rect 23624 13484 24409 13512
rect 23624 13472 23630 13484
rect 24397 13481 24409 13484
rect 24443 13481 24455 13515
rect 24397 13475 24455 13481
rect 21818 13404 21824 13456
rect 21876 13444 21882 13456
rect 24765 13447 24823 13453
rect 21876 13416 22876 13444
rect 21876 13404 21882 13416
rect 21913 13379 21971 13385
rect 21232 13348 21772 13376
rect 21232 13336 21238 13348
rect 19429 13311 19487 13317
rect 19429 13308 19441 13311
rect 18472 13280 19441 13308
rect 18472 13268 18478 13280
rect 19429 13277 19441 13280
rect 19475 13277 19487 13311
rect 19429 13271 19487 13277
rect 19610 13268 19616 13320
rect 19668 13268 19674 13320
rect 19702 13268 19708 13320
rect 19760 13268 19766 13320
rect 21744 13317 21772 13348
rect 21913 13345 21925 13379
rect 21959 13376 21971 13379
rect 22738 13376 22744 13388
rect 21959 13348 22744 13376
rect 21959 13345 21971 13348
rect 21913 13339 21971 13345
rect 22738 13336 22744 13348
rect 22796 13336 22802 13388
rect 21545 13311 21603 13317
rect 21545 13277 21557 13311
rect 21591 13277 21603 13311
rect 21545 13271 21603 13277
rect 21729 13311 21787 13317
rect 21729 13277 21741 13311
rect 21775 13277 21787 13311
rect 21729 13271 21787 13277
rect 22005 13311 22063 13317
rect 22005 13277 22017 13311
rect 22051 13277 22063 13311
rect 22005 13271 22063 13277
rect 18690 13240 18696 13252
rect 16684 13212 18696 13240
rect 16485 13203 16543 13209
rect 18690 13200 18696 13212
rect 18748 13200 18754 13252
rect 19521 13243 19579 13249
rect 19521 13209 19533 13243
rect 19567 13240 19579 13243
rect 19981 13243 20039 13249
rect 19981 13240 19993 13243
rect 19567 13212 19993 13240
rect 19567 13209 19579 13212
rect 19521 13203 19579 13209
rect 19981 13209 19993 13212
rect 20027 13209 20039 13243
rect 21358 13240 21364 13252
rect 21206 13212 21364 13240
rect 19981 13203 20039 13209
rect 21358 13200 21364 13212
rect 21416 13200 21422 13252
rect 21560 13240 21588 13271
rect 21910 13240 21916 13252
rect 21560 13212 21916 13240
rect 21910 13200 21916 13212
rect 21968 13200 21974 13252
rect 22020 13240 22048 13271
rect 22094 13268 22100 13320
rect 22152 13268 22158 13320
rect 22186 13268 22192 13320
rect 22244 13268 22250 13320
rect 22848 13317 22876 13416
rect 24765 13413 24777 13447
rect 24811 13444 24823 13447
rect 24946 13444 24952 13456
rect 24811 13416 24952 13444
rect 24811 13413 24823 13416
rect 24765 13407 24823 13413
rect 24946 13404 24952 13416
rect 25004 13404 25010 13456
rect 22922 13336 22928 13388
rect 22980 13336 22986 13388
rect 23198 13336 23204 13388
rect 23256 13336 23262 13388
rect 22833 13311 22891 13317
rect 22833 13277 22845 13311
rect 22879 13277 22891 13311
rect 22833 13271 22891 13277
rect 24210 13268 24216 13320
rect 24268 13308 24274 13320
rect 24578 13308 24584 13320
rect 24268 13280 24584 13308
rect 24268 13268 24274 13280
rect 24578 13268 24584 13280
rect 24636 13268 24642 13320
rect 24673 13311 24731 13317
rect 24673 13277 24685 13311
rect 24719 13277 24731 13311
rect 24673 13271 24731 13277
rect 22278 13240 22284 13252
rect 22020 13212 22284 13240
rect 22278 13200 22284 13212
rect 22336 13200 22342 13252
rect 22554 13200 22560 13252
rect 22612 13240 22618 13252
rect 24026 13240 24032 13252
rect 22612 13212 24032 13240
rect 22612 13200 22618 13212
rect 24026 13200 24032 13212
rect 24084 13200 24090 13252
rect 24688 13240 24716 13271
rect 24762 13268 24768 13320
rect 24820 13308 24826 13320
rect 24857 13311 24915 13317
rect 24857 13308 24869 13311
rect 24820 13280 24869 13308
rect 24820 13268 24826 13280
rect 24857 13277 24869 13280
rect 24903 13277 24915 13311
rect 24857 13271 24915 13277
rect 24669 13212 24716 13240
rect 15212 13144 15516 13172
rect 16022 13132 16028 13184
rect 16080 13172 16086 13184
rect 20254 13172 20260 13184
rect 16080 13144 20260 13172
rect 16080 13132 16086 13144
rect 20254 13132 20260 13144
rect 20312 13132 20318 13184
rect 21634 13132 21640 13184
rect 21692 13172 21698 13184
rect 23750 13172 23756 13184
rect 21692 13144 23756 13172
rect 21692 13132 21698 13144
rect 23750 13132 23756 13144
rect 23808 13172 23814 13184
rect 24669 13172 24697 13212
rect 23808 13144 24697 13172
rect 23808 13132 23814 13144
rect 1104 13082 28152 13104
rect 1104 13030 4874 13082
rect 4926 13030 4938 13082
rect 4990 13030 5002 13082
rect 5054 13030 5066 13082
rect 5118 13030 5130 13082
rect 5182 13030 28152 13082
rect 1104 13008 28152 13030
rect 2222 12928 2228 12980
rect 2280 12928 2286 12980
rect 5258 12928 5264 12980
rect 5316 12968 5322 12980
rect 6549 12971 6607 12977
rect 5316 12940 5396 12968
rect 5316 12928 5322 12940
rect 5368 12900 5396 12940
rect 6549 12937 6561 12971
rect 6595 12968 6607 12971
rect 7098 12968 7104 12980
rect 6595 12940 7104 12968
rect 6595 12937 6607 12940
rect 6549 12931 6607 12937
rect 7098 12928 7104 12940
rect 7156 12928 7162 12980
rect 7285 12971 7343 12977
rect 7285 12937 7297 12971
rect 7331 12968 7343 12971
rect 8294 12968 8300 12980
rect 7331 12940 8300 12968
rect 7331 12937 7343 12940
rect 7285 12931 7343 12937
rect 8294 12928 8300 12940
rect 8352 12928 8358 12980
rect 12710 12928 12716 12980
rect 12768 12968 12774 12980
rect 13189 12971 13247 12977
rect 13189 12968 13201 12971
rect 12768 12940 13201 12968
rect 12768 12928 12774 12940
rect 13189 12937 13201 12940
rect 13235 12937 13247 12971
rect 13189 12931 13247 12937
rect 13357 12971 13415 12977
rect 13357 12937 13369 12971
rect 13403 12968 13415 12971
rect 15749 12971 15807 12977
rect 13403 12940 14964 12968
rect 13403 12937 13415 12940
rect 13357 12931 13415 12937
rect 14936 12912 14964 12940
rect 15749 12937 15761 12971
rect 15795 12968 15807 12971
rect 16390 12968 16396 12980
rect 15795 12940 16396 12968
rect 15795 12937 15807 12940
rect 15749 12931 15807 12937
rect 16390 12928 16396 12940
rect 16448 12928 16454 12980
rect 17770 12928 17776 12980
rect 17828 12968 17834 12980
rect 18690 12968 18696 12980
rect 17828 12940 18696 12968
rect 17828 12928 17834 12940
rect 18690 12928 18696 12940
rect 18748 12928 18754 12980
rect 20162 12968 20168 12980
rect 19812 12940 20168 12968
rect 19812 12912 19840 12940
rect 20162 12928 20168 12940
rect 20220 12928 20226 12980
rect 22189 12971 22247 12977
rect 22189 12937 22201 12971
rect 22235 12968 22247 12971
rect 22370 12968 22376 12980
rect 22235 12940 22376 12968
rect 22235 12937 22247 12940
rect 22189 12931 22247 12937
rect 22370 12928 22376 12940
rect 22428 12928 22434 12980
rect 22738 12928 22744 12980
rect 22796 12968 22802 12980
rect 24854 12968 24860 12980
rect 22796 12940 24860 12968
rect 22796 12928 22802 12940
rect 5368 12872 6408 12900
rect 2130 12792 2136 12844
rect 2188 12832 2194 12844
rect 2225 12835 2283 12841
rect 2225 12832 2237 12835
rect 2188 12804 2237 12832
rect 2188 12792 2194 12804
rect 2225 12801 2237 12804
rect 2271 12801 2283 12835
rect 2225 12795 2283 12801
rect 2406 12792 2412 12844
rect 2464 12792 2470 12844
rect 4706 12792 4712 12844
rect 4764 12832 4770 12844
rect 5169 12835 5227 12841
rect 5169 12832 5181 12835
rect 4764 12804 5181 12832
rect 4764 12792 4770 12804
rect 5169 12801 5181 12804
rect 5215 12801 5227 12835
rect 5368 12818 5396 12872
rect 6380 12841 6408 12872
rect 12986 12860 12992 12912
rect 13044 12860 13050 12912
rect 14918 12860 14924 12912
rect 14976 12900 14982 12912
rect 14976 12872 15608 12900
rect 14976 12860 14982 12872
rect 6365 12835 6423 12841
rect 5169 12795 5227 12801
rect 6365 12801 6377 12835
rect 6411 12801 6423 12835
rect 6365 12795 6423 12801
rect 6549 12835 6607 12841
rect 6549 12801 6561 12835
rect 6595 12801 6607 12835
rect 6549 12795 6607 12801
rect 5184 12696 5212 12795
rect 6178 12724 6184 12776
rect 6236 12724 6242 12776
rect 6564 12696 6592 12795
rect 7190 12792 7196 12844
rect 7248 12792 7254 12844
rect 7377 12835 7435 12841
rect 7377 12801 7389 12835
rect 7423 12832 7435 12835
rect 7466 12832 7472 12844
rect 7423 12804 7472 12832
rect 7423 12801 7435 12804
rect 7377 12795 7435 12801
rect 7466 12792 7472 12804
rect 7524 12832 7530 12844
rect 7524 12804 7682 12832
rect 7524 12792 7530 12804
rect 8478 12792 8484 12844
rect 8536 12832 8542 12844
rect 8573 12835 8631 12841
rect 8573 12832 8585 12835
rect 8536 12804 8585 12832
rect 8536 12792 8542 12804
rect 8573 12801 8585 12804
rect 8619 12832 8631 12835
rect 9401 12835 9459 12841
rect 9401 12832 9413 12835
rect 8619 12804 9413 12832
rect 8619 12801 8631 12804
rect 8573 12795 8631 12801
rect 9401 12801 9413 12804
rect 9447 12832 9459 12835
rect 9582 12832 9588 12844
rect 9447 12804 9588 12832
rect 9447 12801 9459 12804
rect 9401 12795 9459 12801
rect 9582 12792 9588 12804
rect 9640 12792 9646 12844
rect 13004 12832 13032 12860
rect 15580 12844 15608 12872
rect 15838 12860 15844 12912
rect 15896 12900 15902 12912
rect 19794 12900 19800 12912
rect 15896 12872 19800 12900
rect 15896 12860 15902 12872
rect 19794 12860 19800 12872
rect 19852 12860 19858 12912
rect 20070 12860 20076 12912
rect 20128 12860 20134 12912
rect 21634 12900 21640 12912
rect 20180 12872 21640 12900
rect 13538 12832 13544 12844
rect 13004 12804 13544 12832
rect 13538 12792 13544 12804
rect 13596 12792 13602 12844
rect 14642 12792 14648 12844
rect 14700 12832 14706 12844
rect 15105 12835 15163 12841
rect 15105 12832 15117 12835
rect 14700 12804 15117 12832
rect 14700 12792 14706 12804
rect 15105 12801 15117 12804
rect 15151 12832 15163 12835
rect 15378 12832 15384 12844
rect 15151 12804 15384 12832
rect 15151 12801 15163 12804
rect 15105 12795 15163 12801
rect 15378 12792 15384 12804
rect 15436 12792 15442 12844
rect 15562 12792 15568 12844
rect 15620 12792 15626 12844
rect 16025 12835 16083 12841
rect 16025 12801 16037 12835
rect 16071 12832 16083 12835
rect 16114 12832 16120 12844
rect 16071 12804 16120 12832
rect 16071 12801 16083 12804
rect 16025 12795 16083 12801
rect 16114 12792 16120 12804
rect 16172 12792 16178 12844
rect 17313 12835 17371 12841
rect 17313 12801 17325 12835
rect 17359 12832 17371 12835
rect 18506 12832 18512 12844
rect 17359 12804 18512 12832
rect 17359 12801 17371 12804
rect 17313 12795 17371 12801
rect 18506 12792 18512 12804
rect 18564 12792 18570 12844
rect 18785 12835 18843 12841
rect 18785 12801 18797 12835
rect 18831 12832 18843 12835
rect 19610 12832 19616 12844
rect 18831 12804 19616 12832
rect 18831 12801 18843 12804
rect 18785 12795 18843 12801
rect 7208 12764 7236 12792
rect 7745 12767 7803 12773
rect 7745 12764 7757 12767
rect 7208 12736 7757 12764
rect 7745 12733 7757 12736
rect 7791 12733 7803 12767
rect 7745 12727 7803 12733
rect 9493 12767 9551 12773
rect 9493 12733 9505 12767
rect 9539 12764 9551 12767
rect 9674 12764 9680 12776
rect 9539 12736 9680 12764
rect 9539 12733 9551 12736
rect 9493 12727 9551 12733
rect 9674 12724 9680 12736
rect 9732 12724 9738 12776
rect 10045 12767 10103 12773
rect 10045 12733 10057 12767
rect 10091 12764 10103 12767
rect 10962 12764 10968 12776
rect 10091 12736 10968 12764
rect 10091 12733 10103 12736
rect 10045 12727 10103 12733
rect 10962 12724 10968 12736
rect 11020 12724 11026 12776
rect 18800 12764 18828 12795
rect 19610 12792 19616 12804
rect 19668 12792 19674 12844
rect 19702 12792 19708 12844
rect 19760 12792 19766 12844
rect 20180 12764 20208 12872
rect 21634 12860 21640 12872
rect 21692 12860 21698 12912
rect 22278 12860 22284 12912
rect 22336 12900 22342 12912
rect 22336 12872 22600 12900
rect 22336 12860 22342 12872
rect 20346 12792 20352 12844
rect 20404 12832 20410 12844
rect 20530 12832 20536 12844
rect 20404 12804 20536 12832
rect 20404 12792 20410 12804
rect 20530 12792 20536 12804
rect 20588 12792 20594 12844
rect 20717 12835 20775 12841
rect 20717 12801 20729 12835
rect 20763 12832 20775 12835
rect 20806 12832 20812 12844
rect 20763 12804 20812 12832
rect 20763 12801 20775 12804
rect 20717 12795 20775 12801
rect 15764 12736 18828 12764
rect 18892 12736 20208 12764
rect 5184 12668 6592 12696
rect 10980 12696 11008 12724
rect 15764 12696 15792 12736
rect 10980 12668 15792 12696
rect 15838 12656 15844 12708
rect 15896 12696 15902 12708
rect 16209 12699 16267 12705
rect 16209 12696 16221 12699
rect 15896 12668 16221 12696
rect 15896 12656 15902 12668
rect 16209 12665 16221 12668
rect 16255 12696 16267 12699
rect 18892 12696 18920 12736
rect 20254 12724 20260 12776
rect 20312 12764 20318 12776
rect 20732 12764 20760 12795
rect 20806 12792 20812 12804
rect 20864 12792 20870 12844
rect 20901 12835 20959 12841
rect 20901 12801 20913 12835
rect 20947 12801 20959 12835
rect 20901 12795 20959 12801
rect 20312 12736 20760 12764
rect 20916 12764 20944 12795
rect 20990 12792 20996 12844
rect 21048 12792 21054 12844
rect 21174 12792 21180 12844
rect 21232 12832 21238 12844
rect 21821 12835 21879 12841
rect 21821 12832 21833 12835
rect 21232 12804 21833 12832
rect 21232 12792 21238 12804
rect 21821 12801 21833 12804
rect 21867 12801 21879 12835
rect 21821 12795 21879 12801
rect 22002 12792 22008 12844
rect 22060 12792 22066 12844
rect 22465 12835 22523 12841
rect 22465 12801 22477 12835
rect 22511 12801 22523 12835
rect 22572 12832 22600 12872
rect 22830 12860 22836 12912
rect 22888 12900 22894 12912
rect 22925 12903 22983 12909
rect 22925 12900 22937 12903
rect 22888 12872 22937 12900
rect 22888 12860 22894 12872
rect 22925 12869 22937 12872
rect 22971 12869 22983 12903
rect 22925 12863 22983 12869
rect 23308 12872 23888 12900
rect 23308 12832 23336 12872
rect 22572 12804 23336 12832
rect 22465 12795 22523 12801
rect 21192 12764 21220 12792
rect 20916 12736 21220 12764
rect 20312 12724 20318 12736
rect 22094 12724 22100 12776
rect 22152 12764 22158 12776
rect 22281 12767 22339 12773
rect 22281 12764 22293 12767
rect 22152 12736 22293 12764
rect 22152 12724 22158 12736
rect 22281 12733 22293 12736
rect 22327 12733 22339 12767
rect 22281 12727 22339 12733
rect 22186 12696 22192 12708
rect 16255 12668 18920 12696
rect 20353 12668 22192 12696
rect 16255 12665 16267 12668
rect 16209 12659 16267 12665
rect 12802 12588 12808 12640
rect 12860 12628 12866 12640
rect 13173 12631 13231 12637
rect 13173 12628 13185 12631
rect 12860 12600 13185 12628
rect 12860 12588 12866 12600
rect 13173 12597 13185 12600
rect 13219 12628 13231 12631
rect 13262 12628 13268 12640
rect 13219 12600 13268 12628
rect 13219 12597 13231 12600
rect 13173 12591 13231 12597
rect 13262 12588 13268 12600
rect 13320 12588 13326 12640
rect 15197 12631 15255 12637
rect 15197 12597 15209 12631
rect 15243 12628 15255 12631
rect 15286 12628 15292 12640
rect 15243 12600 15292 12628
rect 15243 12597 15255 12600
rect 15197 12591 15255 12597
rect 15286 12588 15292 12600
rect 15344 12628 15350 12640
rect 15654 12628 15660 12640
rect 15344 12600 15660 12628
rect 15344 12588 15350 12600
rect 15654 12588 15660 12600
rect 15712 12588 15718 12640
rect 17034 12588 17040 12640
rect 17092 12588 17098 12640
rect 19518 12588 19524 12640
rect 19576 12628 19582 12640
rect 19886 12628 19892 12640
rect 19576 12600 19892 12628
rect 19576 12588 19582 12600
rect 19886 12588 19892 12600
rect 19944 12588 19950 12640
rect 20073 12631 20131 12637
rect 20073 12597 20085 12631
rect 20119 12628 20131 12631
rect 20162 12628 20168 12640
rect 20119 12600 20168 12628
rect 20119 12597 20131 12600
rect 20073 12591 20131 12597
rect 20162 12588 20168 12600
rect 20220 12588 20226 12640
rect 20257 12631 20315 12637
rect 20257 12597 20269 12631
rect 20303 12628 20315 12631
rect 20353 12628 20381 12668
rect 22186 12656 22192 12668
rect 22244 12696 22250 12708
rect 22480 12696 22508 12795
rect 23382 12792 23388 12844
rect 23440 12792 23446 12844
rect 23860 12841 23888 12872
rect 24026 12860 24032 12912
rect 24084 12900 24090 12912
rect 24121 12903 24179 12909
rect 24121 12900 24133 12903
rect 24084 12872 24133 12900
rect 24084 12860 24090 12872
rect 24121 12869 24133 12872
rect 24167 12869 24179 12903
rect 24121 12863 24179 12869
rect 24228 12841 24256 12940
rect 24854 12928 24860 12940
rect 24912 12928 24918 12980
rect 23845 12835 23903 12841
rect 23845 12801 23857 12835
rect 23891 12801 23903 12835
rect 23845 12795 23903 12801
rect 24213 12835 24271 12841
rect 24213 12801 24225 12835
rect 24259 12801 24271 12835
rect 24213 12795 24271 12801
rect 23293 12767 23351 12773
rect 23293 12733 23305 12767
rect 23339 12764 23351 12767
rect 23566 12764 23572 12776
rect 23339 12736 23572 12764
rect 23339 12733 23351 12736
rect 23293 12727 23351 12733
rect 23566 12724 23572 12736
rect 23624 12724 23630 12776
rect 23661 12767 23719 12773
rect 23661 12733 23673 12767
rect 23707 12733 23719 12767
rect 23661 12727 23719 12733
rect 22244 12668 22508 12696
rect 22649 12699 22707 12705
rect 22244 12656 22250 12668
rect 22649 12665 22661 12699
rect 22695 12696 22707 12699
rect 23676 12696 23704 12727
rect 22695 12668 23704 12696
rect 22695 12665 22707 12668
rect 22649 12659 22707 12665
rect 20303 12600 20381 12628
rect 20303 12597 20315 12600
rect 20257 12591 20315 12597
rect 20714 12588 20720 12640
rect 20772 12588 20778 12640
rect 21082 12588 21088 12640
rect 21140 12588 21146 12640
rect 23198 12588 23204 12640
rect 23256 12588 23262 12640
rect 23290 12588 23296 12640
rect 23348 12628 23354 12640
rect 23569 12631 23627 12637
rect 23569 12628 23581 12631
rect 23348 12600 23581 12628
rect 23348 12588 23354 12600
rect 23569 12597 23581 12600
rect 23615 12597 23627 12631
rect 23676 12628 23704 12668
rect 24302 12628 24308 12640
rect 23676 12600 24308 12628
rect 23569 12591 23627 12597
rect 24302 12588 24308 12600
rect 24360 12588 24366 12640
rect 1104 12538 28152 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 28152 12538
rect 1104 12464 28152 12486
rect 11146 12384 11152 12436
rect 11204 12424 11210 12436
rect 12345 12427 12403 12433
rect 12345 12424 12357 12427
rect 11204 12396 12357 12424
rect 11204 12384 11210 12396
rect 12345 12393 12357 12396
rect 12391 12393 12403 12427
rect 12345 12387 12403 12393
rect 15378 12384 15384 12436
rect 15436 12424 15442 12436
rect 15565 12427 15623 12433
rect 15565 12424 15577 12427
rect 15436 12396 15577 12424
rect 15436 12384 15442 12396
rect 15565 12393 15577 12396
rect 15611 12393 15623 12427
rect 15838 12424 15844 12436
rect 15565 12387 15623 12393
rect 15672 12396 15844 12424
rect 1854 12316 1860 12368
rect 1912 12356 1918 12368
rect 2682 12356 2688 12368
rect 1912 12328 2688 12356
rect 1912 12316 1918 12328
rect 1964 12297 1992 12328
rect 2682 12316 2688 12328
rect 2740 12316 2746 12368
rect 13722 12316 13728 12368
rect 13780 12356 13786 12368
rect 15672 12356 15700 12396
rect 15838 12384 15844 12396
rect 15896 12384 15902 12436
rect 15930 12384 15936 12436
rect 15988 12424 15994 12436
rect 19245 12427 19303 12433
rect 15988 12396 16160 12424
rect 15988 12384 15994 12396
rect 13780 12328 15700 12356
rect 15749 12359 15807 12365
rect 13780 12316 13786 12328
rect 15749 12325 15761 12359
rect 15795 12356 15807 12359
rect 15795 12328 16068 12356
rect 15795 12325 15807 12328
rect 15749 12319 15807 12325
rect 1949 12291 2007 12297
rect 1949 12257 1961 12291
rect 1995 12257 2007 12291
rect 1949 12251 2007 12257
rect 2225 12291 2283 12297
rect 2225 12257 2237 12291
rect 2271 12288 2283 12291
rect 2406 12288 2412 12300
rect 2271 12260 2412 12288
rect 2271 12257 2283 12260
rect 2225 12251 2283 12257
rect 2406 12248 2412 12260
rect 2464 12248 2470 12300
rect 6178 12248 6184 12300
rect 6236 12288 6242 12300
rect 6549 12291 6607 12297
rect 6549 12288 6561 12291
rect 6236 12260 6561 12288
rect 6236 12248 6242 12260
rect 6549 12257 6561 12260
rect 6595 12257 6607 12291
rect 6549 12251 6607 12257
rect 7466 12248 7472 12300
rect 7524 12248 7530 12300
rect 12713 12291 12771 12297
rect 12713 12257 12725 12291
rect 12759 12288 12771 12291
rect 12894 12288 12900 12300
rect 12759 12260 12900 12288
rect 12759 12257 12771 12260
rect 12713 12251 12771 12257
rect 12894 12248 12900 12260
rect 12952 12248 12958 12300
rect 14090 12248 14096 12300
rect 14148 12288 14154 12300
rect 15838 12288 15844 12300
rect 14148 12260 15844 12288
rect 14148 12248 14154 12260
rect 15838 12248 15844 12260
rect 15896 12248 15902 12300
rect 16040 12297 16068 12328
rect 16025 12291 16083 12297
rect 16025 12257 16037 12291
rect 16071 12257 16083 12291
rect 16025 12251 16083 12257
rect 16132 12288 16160 12396
rect 19245 12393 19257 12427
rect 19291 12424 19303 12427
rect 19426 12424 19432 12436
rect 19291 12396 19432 12424
rect 19291 12393 19303 12396
rect 19245 12387 19303 12393
rect 19426 12384 19432 12396
rect 19484 12384 19490 12436
rect 16574 12316 16580 12368
rect 16632 12356 16638 12368
rect 17678 12356 17684 12368
rect 16632 12328 17684 12356
rect 16632 12316 16638 12328
rect 17678 12316 17684 12328
rect 17736 12316 17742 12368
rect 18690 12316 18696 12368
rect 18748 12356 18754 12368
rect 19613 12359 19671 12365
rect 19613 12356 19625 12359
rect 18748 12328 19625 12356
rect 18748 12316 18754 12328
rect 19613 12325 19625 12328
rect 19659 12325 19671 12359
rect 19613 12319 19671 12325
rect 16850 12288 16856 12300
rect 16132 12260 16856 12288
rect 1857 12223 1915 12229
rect 1857 12189 1869 12223
rect 1903 12220 1915 12223
rect 2038 12220 2044 12232
rect 1903 12192 2044 12220
rect 1903 12189 1915 12192
rect 1857 12183 1915 12189
rect 2038 12180 2044 12192
rect 2096 12180 2102 12232
rect 2130 12180 2136 12232
rect 2188 12220 2194 12232
rect 2501 12223 2559 12229
rect 2501 12220 2513 12223
rect 2188 12192 2513 12220
rect 2188 12180 2194 12192
rect 2501 12189 2513 12192
rect 2547 12189 2559 12223
rect 2501 12183 2559 12189
rect 6095 12223 6153 12229
rect 6095 12189 6107 12223
rect 6141 12220 6153 12223
rect 6196 12220 6224 12248
rect 6141 12192 6224 12220
rect 6273 12223 6331 12229
rect 6141 12189 6153 12192
rect 6095 12183 6153 12189
rect 6273 12189 6285 12223
rect 6319 12220 6331 12223
rect 6641 12223 6699 12229
rect 6641 12220 6653 12223
rect 6319 12192 6653 12220
rect 6319 12189 6331 12192
rect 6273 12183 6331 12189
rect 6641 12189 6653 12192
rect 6687 12220 6699 12223
rect 8478 12220 8484 12232
rect 6687 12192 8484 12220
rect 6687 12189 6699 12192
rect 6641 12183 6699 12189
rect 8478 12180 8484 12192
rect 8536 12180 8542 12232
rect 12526 12180 12532 12232
rect 12584 12180 12590 12232
rect 12618 12180 12624 12232
rect 12676 12180 12682 12232
rect 12805 12223 12863 12229
rect 12805 12189 12817 12223
rect 12851 12220 12863 12223
rect 13170 12220 13176 12232
rect 12851 12192 13176 12220
rect 12851 12189 12863 12192
rect 12805 12183 12863 12189
rect 13170 12180 13176 12192
rect 13228 12180 13234 12232
rect 12710 12112 12716 12164
rect 12768 12152 12774 12164
rect 14108 12152 14136 12248
rect 16132 12229 16160 12260
rect 16850 12248 16856 12260
rect 16908 12248 16914 12300
rect 19521 12291 19579 12297
rect 19521 12257 19533 12291
rect 19567 12288 19579 12291
rect 20714 12288 20720 12300
rect 19567 12260 20720 12288
rect 19567 12257 19579 12260
rect 19521 12251 19579 12257
rect 20714 12248 20720 12260
rect 20772 12248 20778 12300
rect 16117 12223 16175 12229
rect 15396 12192 16068 12220
rect 15396 12164 15424 12192
rect 12768 12124 14136 12152
rect 12768 12112 12774 12124
rect 15378 12112 15384 12164
rect 15436 12112 15442 12164
rect 15562 12112 15568 12164
rect 15620 12161 15626 12164
rect 15620 12155 15639 12161
rect 15627 12121 15639 12155
rect 15620 12115 15639 12121
rect 15620 12112 15626 12115
rect 15838 12112 15844 12164
rect 15896 12112 15902 12164
rect 16040 12152 16068 12192
rect 16117 12189 16129 12223
rect 16163 12189 16175 12223
rect 16117 12183 16175 12189
rect 16482 12180 16488 12232
rect 16540 12220 16546 12232
rect 17037 12223 17095 12229
rect 17037 12220 17049 12223
rect 16540 12192 17049 12220
rect 16540 12180 16546 12192
rect 17037 12189 17049 12192
rect 17083 12189 17095 12223
rect 17037 12183 17095 12189
rect 18785 12223 18843 12229
rect 18785 12189 18797 12223
rect 18831 12220 18843 12223
rect 19334 12220 19340 12232
rect 18831 12192 19340 12220
rect 18831 12189 18843 12192
rect 18785 12183 18843 12189
rect 19334 12180 19340 12192
rect 19392 12180 19398 12232
rect 19429 12223 19487 12229
rect 19429 12189 19441 12223
rect 19475 12189 19487 12223
rect 19429 12183 19487 12189
rect 19705 12223 19763 12229
rect 19705 12189 19717 12223
rect 19751 12220 19763 12223
rect 19794 12220 19800 12232
rect 19751 12192 19800 12220
rect 19751 12189 19763 12192
rect 19705 12183 19763 12189
rect 16574 12152 16580 12164
rect 16040 12124 16580 12152
rect 16574 12112 16580 12124
rect 16632 12112 16638 12164
rect 16761 12155 16819 12161
rect 16761 12121 16773 12155
rect 16807 12152 16819 12155
rect 16942 12152 16948 12164
rect 16807 12124 16948 12152
rect 16807 12121 16819 12124
rect 16761 12115 16819 12121
rect 16942 12112 16948 12124
rect 17000 12112 17006 12164
rect 2866 12044 2872 12096
rect 2924 12044 2930 12096
rect 6273 12087 6331 12093
rect 6273 12053 6285 12087
rect 6319 12084 6331 12087
rect 7006 12084 7012 12096
rect 6319 12056 7012 12084
rect 6319 12053 6331 12056
rect 6273 12047 6331 12053
rect 7006 12044 7012 12056
rect 7064 12044 7070 12096
rect 15930 12044 15936 12096
rect 15988 12084 15994 12096
rect 16301 12087 16359 12093
rect 16301 12084 16313 12087
rect 15988 12056 16313 12084
rect 15988 12044 15994 12056
rect 16301 12053 16313 12056
rect 16347 12053 16359 12087
rect 16301 12047 16359 12053
rect 16485 12087 16543 12093
rect 16485 12053 16497 12087
rect 16531 12084 16543 12087
rect 18414 12084 18420 12096
rect 16531 12056 18420 12084
rect 16531 12053 16543 12056
rect 16485 12047 16543 12053
rect 18414 12044 18420 12056
rect 18472 12044 18478 12096
rect 19444 12084 19472 12183
rect 19794 12180 19800 12192
rect 19852 12180 19858 12232
rect 19889 12223 19947 12229
rect 19889 12189 19901 12223
rect 19935 12220 19947 12223
rect 21082 12220 21088 12232
rect 19935 12192 21088 12220
rect 19935 12189 19947 12192
rect 19889 12183 19947 12189
rect 21082 12180 21088 12192
rect 21140 12180 21146 12232
rect 19518 12112 19524 12164
rect 19576 12152 19582 12164
rect 20257 12155 20315 12161
rect 20257 12152 20269 12155
rect 19576 12124 20269 12152
rect 19576 12112 19582 12124
rect 20257 12121 20269 12124
rect 20303 12121 20315 12155
rect 21266 12152 21272 12164
rect 20257 12115 20315 12121
rect 20456 12124 21272 12152
rect 20456 12084 20484 12124
rect 21266 12112 21272 12124
rect 21324 12112 21330 12164
rect 19444 12056 20484 12084
rect 20530 12044 20536 12096
rect 20588 12084 20594 12096
rect 21545 12087 21603 12093
rect 21545 12084 21557 12087
rect 20588 12056 21557 12084
rect 20588 12044 20594 12056
rect 21545 12053 21557 12056
rect 21591 12084 21603 12087
rect 23474 12084 23480 12096
rect 21591 12056 23480 12084
rect 21591 12053 21603 12056
rect 21545 12047 21603 12053
rect 23474 12044 23480 12056
rect 23532 12084 23538 12096
rect 24670 12084 24676 12096
rect 23532 12056 24676 12084
rect 23532 12044 23538 12056
rect 24670 12044 24676 12056
rect 24728 12044 24734 12096
rect 1104 11994 28152 12016
rect 1104 11942 4874 11994
rect 4926 11942 4938 11994
rect 4990 11942 5002 11994
rect 5054 11942 5066 11994
rect 5118 11942 5130 11994
rect 5182 11942 28152 11994
rect 1104 11920 28152 11942
rect 4522 11880 4528 11892
rect 3896 11852 4528 11880
rect 842 11704 848 11756
rect 900 11744 906 11756
rect 3896 11753 3924 11852
rect 4522 11840 4528 11852
rect 4580 11840 4586 11892
rect 9585 11883 9643 11889
rect 9585 11849 9597 11883
rect 9631 11880 9643 11883
rect 12434 11880 12440 11892
rect 9631 11852 12440 11880
rect 9631 11849 9643 11852
rect 9585 11843 9643 11849
rect 12434 11840 12440 11852
rect 12492 11840 12498 11892
rect 12529 11883 12587 11889
rect 12529 11849 12541 11883
rect 12575 11880 12587 11883
rect 12618 11880 12624 11892
rect 12575 11852 12624 11880
rect 12575 11849 12587 11852
rect 12529 11843 12587 11849
rect 12618 11840 12624 11852
rect 12676 11840 12682 11892
rect 12986 11840 12992 11892
rect 13044 11840 13050 11892
rect 13170 11840 13176 11892
rect 13228 11840 13234 11892
rect 13354 11840 13360 11892
rect 13412 11880 13418 11892
rect 13412 11852 14044 11880
rect 13412 11840 13418 11852
rect 4706 11772 4712 11824
rect 4764 11772 4770 11824
rect 4798 11772 4804 11824
rect 4856 11812 4862 11824
rect 4856 11784 5396 11812
rect 4856 11772 4862 11784
rect 4341 11757 4399 11763
rect 4341 11754 4353 11757
rect 1397 11747 1455 11753
rect 1397 11744 1409 11747
rect 900 11716 1409 11744
rect 900 11704 906 11716
rect 1397 11713 1409 11716
rect 1443 11713 1455 11747
rect 1397 11707 1455 11713
rect 3881 11747 3939 11753
rect 3881 11713 3893 11747
rect 3927 11713 3939 11747
rect 3881 11707 3939 11713
rect 4264 11726 4353 11754
rect 1673 11679 1731 11685
rect 1673 11645 1685 11679
rect 1719 11676 1731 11679
rect 1946 11676 1952 11688
rect 1719 11648 1952 11676
rect 1719 11645 1731 11648
rect 1673 11639 1731 11645
rect 1946 11636 1952 11648
rect 2004 11636 2010 11688
rect 3786 11636 3792 11688
rect 3844 11676 3850 11688
rect 4264 11676 4292 11726
rect 4341 11723 4353 11726
rect 4387 11723 4399 11757
rect 5368 11756 5396 11784
rect 7650 11772 7656 11824
rect 7708 11812 7714 11824
rect 8941 11815 8999 11821
rect 8941 11812 8953 11815
rect 7708 11784 8953 11812
rect 7708 11772 7714 11784
rect 4341 11717 4399 11723
rect 4522 11704 4528 11756
rect 4580 11704 4586 11756
rect 4617 11747 4675 11753
rect 4617 11713 4629 11747
rect 4663 11713 4675 11747
rect 4890 11744 4896 11756
rect 4617 11707 4675 11713
rect 4724 11716 4896 11744
rect 3844 11648 4292 11676
rect 4433 11679 4491 11685
rect 3844 11636 3850 11648
rect 4433 11645 4445 11679
rect 4479 11676 4491 11679
rect 4632 11676 4660 11707
rect 4479 11648 4660 11676
rect 4479 11645 4491 11648
rect 4433 11639 4491 11645
rect 4249 11611 4307 11617
rect 4249 11577 4261 11611
rect 4295 11608 4307 11611
rect 4724 11608 4752 11716
rect 4890 11704 4896 11716
rect 4948 11704 4954 11756
rect 5169 11747 5227 11753
rect 5169 11713 5181 11747
rect 5215 11713 5227 11747
rect 5169 11707 5227 11713
rect 5184 11676 5212 11707
rect 5350 11704 5356 11756
rect 5408 11704 5414 11756
rect 8680 11753 8708 11784
rect 8941 11781 8953 11784
rect 8987 11812 8999 11815
rect 8987 11784 9720 11812
rect 8987 11781 8999 11784
rect 8941 11775 8999 11781
rect 8481 11747 8539 11753
rect 8481 11713 8493 11747
rect 8527 11713 8539 11747
rect 8481 11707 8539 11713
rect 8665 11747 8723 11753
rect 8665 11713 8677 11747
rect 8711 11713 8723 11747
rect 8665 11707 8723 11713
rect 5534 11676 5540 11688
rect 5184 11648 5540 11676
rect 5534 11636 5540 11648
rect 5592 11636 5598 11688
rect 4295 11580 4752 11608
rect 8496 11608 8524 11707
rect 8754 11704 8760 11756
rect 8812 11704 8818 11756
rect 9692 11753 9720 11784
rect 10962 11772 10968 11824
rect 11020 11772 11026 11824
rect 11054 11772 11060 11824
rect 11112 11812 11118 11824
rect 11165 11815 11223 11821
rect 11165 11812 11177 11815
rect 11112 11784 11177 11812
rect 11112 11772 11118 11784
rect 11165 11781 11177 11784
rect 11211 11781 11223 11815
rect 11165 11775 11223 11781
rect 9125 11747 9183 11753
rect 9125 11713 9137 11747
rect 9171 11744 9183 11747
rect 9401 11747 9459 11753
rect 9401 11744 9413 11747
rect 9171 11716 9413 11744
rect 9171 11713 9183 11716
rect 9125 11707 9183 11713
rect 9401 11713 9413 11716
rect 9447 11713 9459 11747
rect 9401 11707 9459 11713
rect 9585 11747 9643 11753
rect 9585 11713 9597 11747
rect 9631 11713 9643 11747
rect 9585 11707 9643 11713
rect 9677 11747 9735 11753
rect 9677 11713 9689 11747
rect 9723 11713 9735 11747
rect 9677 11707 9735 11713
rect 8573 11679 8631 11685
rect 8573 11645 8585 11679
rect 8619 11676 8631 11679
rect 9214 11676 9220 11688
rect 8619 11648 9220 11676
rect 8619 11645 8631 11648
rect 8573 11639 8631 11645
rect 9214 11636 9220 11648
rect 9272 11676 9278 11688
rect 9600 11676 9628 11707
rect 9858 11704 9864 11756
rect 9916 11744 9922 11756
rect 10226 11744 10232 11756
rect 9916 11716 10232 11744
rect 9916 11704 9922 11716
rect 10226 11704 10232 11716
rect 10284 11704 10290 11756
rect 12250 11704 12256 11756
rect 12308 11744 12314 11756
rect 13004 11753 13032 11840
rect 13906 11812 13912 11824
rect 13096 11784 13492 11812
rect 13096 11756 13124 11784
rect 12713 11747 12771 11753
rect 12713 11744 12725 11747
rect 12308 11716 12725 11744
rect 12308 11704 12314 11716
rect 12713 11713 12725 11716
rect 12759 11713 12771 11747
rect 12713 11707 12771 11713
rect 12805 11747 12863 11753
rect 12805 11713 12817 11747
rect 12851 11713 12863 11747
rect 12805 11707 12863 11713
rect 12989 11747 13047 11753
rect 12989 11713 13001 11747
rect 13035 11713 13047 11747
rect 12989 11707 13047 11713
rect 9272 11648 9628 11676
rect 9272 11636 9278 11648
rect 9766 11636 9772 11688
rect 9824 11676 9830 11688
rect 9824 11648 12434 11676
rect 9824 11636 9830 11648
rect 8754 11608 8760 11620
rect 8496 11580 8760 11608
rect 4295 11577 4307 11580
rect 4249 11571 4307 11577
rect 8754 11568 8760 11580
rect 8812 11568 8818 11620
rect 11330 11568 11336 11620
rect 11388 11568 11394 11620
rect 12406 11608 12434 11648
rect 12618 11636 12624 11688
rect 12676 11676 12682 11688
rect 12820 11676 12848 11707
rect 13078 11704 13084 11756
rect 13136 11704 13142 11756
rect 13170 11704 13176 11756
rect 13228 11744 13234 11756
rect 13357 11747 13415 11753
rect 13357 11744 13369 11747
rect 13228 11716 13369 11744
rect 13228 11704 13234 11716
rect 13357 11713 13369 11716
rect 13403 11713 13415 11747
rect 13464 11744 13492 11784
rect 13648 11784 13912 11812
rect 13648 11753 13676 11784
rect 13906 11772 13912 11784
rect 13964 11772 13970 11824
rect 14016 11821 14044 11852
rect 14642 11840 14648 11892
rect 14700 11840 14706 11892
rect 15470 11880 15476 11892
rect 15212 11852 15476 11880
rect 14001 11815 14059 11821
rect 14001 11781 14013 11815
rect 14047 11781 14059 11815
rect 14001 11775 14059 11781
rect 14093 11815 14151 11821
rect 14093 11781 14105 11815
rect 14139 11812 14151 11815
rect 14660 11812 14688 11840
rect 14139 11784 14688 11812
rect 14139 11781 14151 11784
rect 14093 11775 14151 11781
rect 13541 11747 13599 11753
rect 13541 11744 13553 11747
rect 13464 11716 13553 11744
rect 13357 11707 13415 11713
rect 13541 11713 13553 11716
rect 13587 11713 13599 11747
rect 13541 11707 13599 11713
rect 13633 11747 13691 11753
rect 13633 11713 13645 11747
rect 13679 11713 13691 11747
rect 13633 11707 13691 11713
rect 13814 11704 13820 11756
rect 13872 11704 13878 11756
rect 12676 11648 12848 11676
rect 12676 11636 12682 11648
rect 13722 11636 13728 11688
rect 13780 11676 13786 11688
rect 14016 11676 14044 11775
rect 14185 11747 14243 11753
rect 14185 11744 14197 11747
rect 13780 11648 14044 11676
rect 14108 11716 14197 11744
rect 13780 11636 13786 11648
rect 14108 11608 14136 11716
rect 14185 11713 14197 11716
rect 14231 11744 14243 11747
rect 14645 11747 14703 11753
rect 14645 11744 14657 11747
rect 14231 11716 14657 11744
rect 14231 11713 14243 11716
rect 14185 11707 14243 11713
rect 14645 11713 14657 11716
rect 14691 11713 14703 11747
rect 14645 11707 14703 11713
rect 12406 11580 14136 11608
rect 15212 11608 15240 11852
rect 15470 11840 15476 11852
rect 15528 11840 15534 11892
rect 15562 11840 15568 11892
rect 15620 11840 15626 11892
rect 19334 11840 19340 11892
rect 19392 11880 19398 11892
rect 19978 11880 19984 11892
rect 19392 11852 19984 11880
rect 19392 11840 19398 11852
rect 19978 11840 19984 11852
rect 20036 11840 20042 11892
rect 20162 11840 20168 11892
rect 20220 11880 20226 11892
rect 20220 11852 23520 11880
rect 20220 11840 20226 11852
rect 16025 11815 16083 11821
rect 15304 11784 15976 11812
rect 15304 11753 15332 11784
rect 15948 11756 15976 11784
rect 16025 11781 16037 11815
rect 16071 11812 16083 11815
rect 18601 11815 18659 11821
rect 18601 11812 18613 11815
rect 16071 11784 18613 11812
rect 16071 11781 16083 11784
rect 16025 11775 16083 11781
rect 18601 11781 18613 11784
rect 18647 11781 18659 11815
rect 18601 11775 18659 11781
rect 19061 11815 19119 11821
rect 19061 11781 19073 11815
rect 19107 11812 19119 11815
rect 22646 11812 22652 11824
rect 19107 11784 22652 11812
rect 19107 11781 19119 11784
rect 19061 11775 19119 11781
rect 15289 11747 15347 11753
rect 15289 11713 15301 11747
rect 15335 11713 15347 11747
rect 15289 11707 15347 11713
rect 15381 11747 15439 11753
rect 15381 11713 15393 11747
rect 15427 11713 15439 11747
rect 15381 11707 15439 11713
rect 15396 11608 15424 11707
rect 15562 11704 15568 11756
rect 15620 11742 15626 11756
rect 15657 11747 15715 11753
rect 15657 11742 15669 11747
rect 15620 11714 15669 11742
rect 15620 11704 15626 11714
rect 15657 11713 15669 11714
rect 15703 11713 15715 11747
rect 15657 11707 15715 11713
rect 15930 11704 15936 11756
rect 15988 11704 15994 11756
rect 15470 11636 15476 11688
rect 15528 11636 15534 11688
rect 16040 11608 16068 11775
rect 22646 11772 22652 11784
rect 22704 11772 22710 11824
rect 23492 11812 23520 11852
rect 23566 11840 23572 11892
rect 23624 11880 23630 11892
rect 23661 11883 23719 11889
rect 23661 11880 23673 11883
rect 23624 11852 23673 11880
rect 23624 11840 23630 11852
rect 23661 11849 23673 11852
rect 23707 11849 23719 11883
rect 25130 11880 25136 11892
rect 23661 11843 23719 11849
rect 23860 11852 25136 11880
rect 23860 11812 23888 11852
rect 25130 11840 25136 11852
rect 25188 11880 25194 11892
rect 25409 11883 25467 11889
rect 25409 11880 25421 11883
rect 25188 11852 25421 11880
rect 25188 11840 25194 11852
rect 25409 11849 25421 11852
rect 25455 11849 25467 11883
rect 25409 11843 25467 11849
rect 23492 11784 23888 11812
rect 23937 11815 23995 11821
rect 23937 11781 23949 11815
rect 23983 11812 23995 11815
rect 24394 11812 24400 11824
rect 23983 11784 24400 11812
rect 23983 11781 23995 11784
rect 23937 11775 23995 11781
rect 24394 11772 24400 11784
rect 24452 11772 24458 11824
rect 16114 11704 16120 11756
rect 16172 11704 16178 11756
rect 16298 11704 16304 11756
rect 16356 11704 16362 11756
rect 16393 11747 16451 11753
rect 16393 11713 16405 11747
rect 16439 11713 16451 11747
rect 16393 11707 16451 11713
rect 15212 11580 15332 11608
rect 15396 11580 16068 11608
rect 9582 11500 9588 11552
rect 9640 11540 9646 11552
rect 9861 11543 9919 11549
rect 9861 11540 9873 11543
rect 9640 11512 9873 11540
rect 9640 11500 9646 11512
rect 9861 11509 9873 11512
rect 9907 11509 9919 11543
rect 9861 11503 9919 11509
rect 11146 11500 11152 11552
rect 11204 11500 11210 11552
rect 13170 11500 13176 11552
rect 13228 11540 13234 11552
rect 13446 11540 13452 11552
rect 13228 11512 13452 11540
rect 13228 11500 13234 11512
rect 13446 11500 13452 11512
rect 13504 11500 13510 11552
rect 13538 11500 13544 11552
rect 13596 11540 13602 11552
rect 13814 11540 13820 11552
rect 13596 11512 13820 11540
rect 13596 11500 13602 11512
rect 13814 11500 13820 11512
rect 13872 11500 13878 11552
rect 14369 11543 14427 11549
rect 14369 11509 14381 11543
rect 14415 11540 14427 11543
rect 14458 11540 14464 11552
rect 14415 11512 14464 11540
rect 14415 11509 14427 11512
rect 14369 11503 14427 11509
rect 14458 11500 14464 11512
rect 14516 11500 14522 11552
rect 14737 11543 14795 11549
rect 14737 11509 14749 11543
rect 14783 11540 14795 11543
rect 15194 11540 15200 11552
rect 14783 11512 15200 11540
rect 14783 11509 14795 11512
rect 14737 11503 14795 11509
rect 15194 11500 15200 11512
rect 15252 11500 15258 11552
rect 15304 11540 15332 11580
rect 15749 11543 15807 11549
rect 15749 11540 15761 11543
rect 15304 11512 15761 11540
rect 15749 11509 15761 11512
rect 15795 11509 15807 11543
rect 15749 11503 15807 11509
rect 16022 11500 16028 11552
rect 16080 11540 16086 11552
rect 16408 11540 16436 11707
rect 16482 11704 16488 11756
rect 16540 11744 16546 11756
rect 17037 11747 17095 11753
rect 17037 11744 17049 11747
rect 16540 11716 17049 11744
rect 16540 11704 16546 11716
rect 17037 11713 17049 11716
rect 17083 11713 17095 11747
rect 17037 11707 17095 11713
rect 17218 11704 17224 11756
rect 17276 11744 17282 11756
rect 18049 11747 18107 11753
rect 18049 11744 18061 11747
rect 17276 11716 18061 11744
rect 17276 11704 17282 11716
rect 18049 11713 18061 11716
rect 18095 11713 18107 11747
rect 18049 11707 18107 11713
rect 18141 11747 18199 11753
rect 18141 11713 18153 11747
rect 18187 11713 18199 11747
rect 18141 11707 18199 11713
rect 18325 11747 18383 11753
rect 18325 11713 18337 11747
rect 18371 11713 18383 11747
rect 18325 11707 18383 11713
rect 18156 11676 18184 11707
rect 17052 11648 18184 11676
rect 18340 11676 18368 11707
rect 18414 11704 18420 11756
rect 18472 11744 18478 11756
rect 19521 11747 19579 11753
rect 18472 11716 18920 11744
rect 18472 11704 18478 11716
rect 18340 11648 18828 11676
rect 17052 11620 17080 11648
rect 17034 11568 17040 11620
rect 17092 11568 17098 11620
rect 16080 11512 16436 11540
rect 16080 11500 16086 11512
rect 16758 11500 16764 11552
rect 16816 11540 16822 11552
rect 16942 11540 16948 11552
rect 16816 11512 16948 11540
rect 16816 11500 16822 11512
rect 16942 11500 16948 11512
rect 17000 11500 17006 11552
rect 18156 11540 18184 11648
rect 18800 11552 18828 11648
rect 18598 11540 18604 11552
rect 18156 11512 18604 11540
rect 18598 11500 18604 11512
rect 18656 11500 18662 11552
rect 18782 11500 18788 11552
rect 18840 11500 18846 11552
rect 18892 11540 18920 11716
rect 19521 11713 19533 11747
rect 19567 11744 19579 11747
rect 20533 11747 20591 11753
rect 19567 11716 20484 11744
rect 19567 11713 19579 11716
rect 19521 11707 19579 11713
rect 19610 11636 19616 11688
rect 19668 11636 19674 11688
rect 20257 11679 20315 11685
rect 20257 11645 20269 11679
rect 20303 11645 20315 11679
rect 20456 11676 20484 11716
rect 20533 11713 20545 11747
rect 20579 11744 20591 11747
rect 21082 11744 21088 11756
rect 20579 11716 21088 11744
rect 20579 11713 20591 11716
rect 20533 11707 20591 11713
rect 21082 11704 21088 11716
rect 21140 11704 21146 11756
rect 23842 11704 23848 11756
rect 23900 11704 23906 11756
rect 24029 11747 24087 11753
rect 24029 11713 24041 11747
rect 24075 11744 24087 11747
rect 24118 11744 24124 11756
rect 24075 11716 24124 11744
rect 24075 11713 24087 11716
rect 24029 11707 24087 11713
rect 24118 11704 24124 11716
rect 24176 11704 24182 11756
rect 24213 11747 24271 11753
rect 24213 11713 24225 11747
rect 24259 11713 24271 11747
rect 24213 11707 24271 11713
rect 20806 11676 20812 11688
rect 20456 11648 20812 11676
rect 20257 11639 20315 11645
rect 19889 11611 19947 11617
rect 19889 11577 19901 11611
rect 19935 11608 19947 11611
rect 19935 11580 20208 11608
rect 19935 11577 19947 11580
rect 19889 11571 19947 11577
rect 19978 11540 19984 11552
rect 18892 11512 19984 11540
rect 19978 11500 19984 11512
rect 20036 11500 20042 11552
rect 20180 11549 20208 11580
rect 20165 11543 20223 11549
rect 20165 11509 20177 11543
rect 20211 11509 20223 11543
rect 20272 11540 20300 11639
rect 20806 11636 20812 11648
rect 20864 11636 20870 11688
rect 24228 11676 24256 11707
rect 24302 11704 24308 11756
rect 24360 11704 24366 11756
rect 24581 11747 24639 11753
rect 24581 11713 24593 11747
rect 24627 11744 24639 11747
rect 24854 11744 24860 11756
rect 24627 11716 24860 11744
rect 24627 11713 24639 11716
rect 24581 11707 24639 11713
rect 24854 11704 24860 11716
rect 24912 11704 24918 11756
rect 25682 11704 25688 11756
rect 25740 11744 25746 11756
rect 26602 11744 26608 11756
rect 25740 11716 26608 11744
rect 25740 11704 25746 11716
rect 26602 11704 26608 11716
rect 26660 11704 26666 11756
rect 24486 11676 24492 11688
rect 24228 11648 24492 11676
rect 24486 11636 24492 11648
rect 24544 11636 24550 11688
rect 20714 11540 20720 11552
rect 20272 11512 20720 11540
rect 20165 11503 20223 11509
rect 20714 11500 20720 11512
rect 20772 11500 20778 11552
rect 24026 11500 24032 11552
rect 24084 11540 24090 11552
rect 24489 11543 24547 11549
rect 24489 11540 24501 11543
rect 24084 11512 24501 11540
rect 24084 11500 24090 11512
rect 24489 11509 24501 11512
rect 24535 11509 24547 11543
rect 24489 11503 24547 11509
rect 1104 11450 28152 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 28152 11450
rect 1104 11376 28152 11398
rect 4341 11339 4399 11345
rect 4341 11305 4353 11339
rect 4387 11336 4399 11339
rect 4614 11336 4620 11348
rect 4387 11308 4620 11336
rect 4387 11305 4399 11308
rect 4341 11299 4399 11305
rect 4614 11296 4620 11308
rect 4672 11296 4678 11348
rect 10321 11339 10379 11345
rect 10321 11305 10333 11339
rect 10367 11336 10379 11339
rect 11054 11336 11060 11348
rect 10367 11308 11060 11336
rect 10367 11305 10379 11308
rect 10321 11299 10379 11305
rect 11054 11296 11060 11308
rect 11112 11296 11118 11348
rect 12158 11296 12164 11348
rect 12216 11296 12222 11348
rect 12526 11296 12532 11348
rect 12584 11336 12590 11348
rect 12713 11339 12771 11345
rect 12713 11336 12725 11339
rect 12584 11308 12725 11336
rect 12584 11296 12590 11308
rect 12713 11305 12725 11308
rect 12759 11305 12771 11339
rect 12713 11299 12771 11305
rect 13170 11296 13176 11348
rect 13228 11336 13234 11348
rect 13630 11336 13636 11348
rect 13228 11308 13636 11336
rect 13228 11296 13234 11308
rect 13630 11296 13636 11308
rect 13688 11296 13694 11348
rect 15565 11339 15623 11345
rect 15565 11305 15577 11339
rect 15611 11336 15623 11339
rect 15838 11336 15844 11348
rect 15611 11308 15844 11336
rect 15611 11305 15623 11308
rect 15565 11299 15623 11305
rect 15838 11296 15844 11308
rect 15896 11296 15902 11348
rect 16390 11336 16396 11348
rect 16040 11308 16396 11336
rect 5445 11271 5503 11277
rect 5445 11268 5457 11271
rect 5000 11240 5457 11268
rect 3053 11203 3111 11209
rect 3053 11169 3065 11203
rect 3099 11200 3111 11203
rect 3881 11203 3939 11209
rect 3881 11200 3893 11203
rect 3099 11172 3893 11200
rect 3099 11169 3111 11172
rect 3053 11163 3111 11169
rect 3881 11169 3893 11172
rect 3927 11169 3939 11203
rect 3881 11163 3939 11169
rect 3973 11203 4031 11209
rect 3973 11169 3985 11203
rect 4019 11200 4031 11203
rect 4798 11200 4804 11212
rect 4019 11172 4804 11200
rect 4019 11169 4031 11172
rect 3973 11163 4031 11169
rect 4798 11160 4804 11172
rect 4856 11160 4862 11212
rect 4890 11160 4896 11212
rect 4948 11160 4954 11212
rect 2866 11092 2872 11144
rect 2924 11132 2930 11144
rect 2961 11135 3019 11141
rect 2961 11132 2973 11135
rect 2924 11104 2973 11132
rect 2924 11092 2930 11104
rect 2961 11101 2973 11104
rect 3007 11101 3019 11135
rect 2961 11095 3019 11101
rect 3142 11092 3148 11144
rect 3200 11092 3206 11144
rect 4065 11135 4123 11141
rect 4065 11101 4077 11135
rect 4111 11101 4123 11135
rect 4065 11095 4123 11101
rect 1946 11024 1952 11076
rect 2004 11064 2010 11076
rect 4080 11064 4108 11095
rect 4154 11092 4160 11144
rect 4212 11092 4218 11144
rect 5000 11141 5028 11240
rect 5445 11237 5457 11240
rect 5491 11237 5503 11271
rect 5445 11231 5503 11237
rect 7190 11228 7196 11280
rect 7248 11228 7254 11280
rect 11422 11228 11428 11280
rect 11480 11268 11486 11280
rect 11480 11240 12204 11268
rect 11480 11228 11486 11240
rect 5350 11160 5356 11212
rect 5408 11200 5414 11212
rect 5408 11172 5672 11200
rect 5408 11160 5414 11172
rect 4985 11135 5043 11141
rect 4985 11101 4997 11135
rect 5031 11101 5043 11135
rect 4985 11095 5043 11101
rect 5445 11135 5503 11141
rect 5445 11101 5457 11135
rect 5491 11132 5503 11135
rect 5534 11132 5540 11144
rect 5491 11104 5540 11132
rect 5491 11101 5503 11104
rect 5445 11095 5503 11101
rect 5534 11092 5540 11104
rect 5592 11092 5598 11144
rect 5644 11141 5672 11172
rect 7558 11160 7564 11212
rect 7616 11160 7622 11212
rect 9309 11203 9367 11209
rect 9309 11169 9321 11203
rect 9355 11200 9367 11203
rect 11606 11200 11612 11212
rect 9355 11172 11612 11200
rect 9355 11169 9367 11172
rect 9309 11163 9367 11169
rect 11606 11160 11612 11172
rect 11664 11160 11670 11212
rect 5629 11135 5687 11141
rect 5629 11101 5641 11135
rect 5675 11101 5687 11135
rect 5629 11095 5687 11101
rect 7469 11135 7527 11141
rect 7469 11101 7481 11135
rect 7515 11132 7527 11135
rect 8570 11132 8576 11144
rect 7515 11104 8576 11132
rect 7515 11101 7527 11104
rect 7469 11095 7527 11101
rect 8570 11092 8576 11104
rect 8628 11092 8634 11144
rect 9493 11135 9551 11141
rect 9493 11101 9505 11135
rect 9539 11132 9551 11135
rect 9582 11132 9588 11144
rect 9539 11104 9588 11132
rect 9539 11101 9551 11104
rect 9493 11095 9551 11101
rect 9582 11092 9588 11104
rect 9640 11092 9646 11144
rect 9677 11135 9735 11141
rect 9677 11101 9689 11135
rect 9723 11132 9735 11135
rect 9766 11132 9772 11144
rect 9723 11104 9772 11132
rect 9723 11101 9735 11104
rect 9677 11095 9735 11101
rect 9766 11092 9772 11104
rect 9824 11132 9830 11144
rect 9950 11132 9956 11144
rect 9824 11104 9956 11132
rect 9824 11092 9830 11104
rect 9950 11092 9956 11104
rect 10008 11092 10014 11144
rect 10594 11092 10600 11144
rect 10652 11132 10658 11144
rect 11514 11132 11520 11144
rect 10652 11104 11520 11132
rect 10652 11092 10658 11104
rect 11514 11092 11520 11104
rect 11572 11092 11578 11144
rect 11808 11141 11836 11240
rect 11882 11160 11888 11212
rect 11940 11200 11946 11212
rect 12176 11200 12204 11240
rect 12894 11228 12900 11280
rect 12952 11268 12958 11280
rect 15470 11268 15476 11280
rect 12952 11240 15476 11268
rect 12952 11228 12958 11240
rect 13648 11212 13676 11240
rect 15470 11228 15476 11240
rect 15528 11268 15534 11280
rect 15930 11268 15936 11280
rect 15528 11240 15936 11268
rect 15528 11228 15534 11240
rect 15930 11228 15936 11240
rect 15988 11228 15994 11280
rect 11940 11172 12112 11200
rect 12176 11172 13032 11200
rect 11940 11160 11946 11172
rect 11793 11135 11851 11141
rect 11793 11101 11805 11135
rect 11839 11101 11851 11135
rect 11793 11095 11851 11101
rect 11974 11092 11980 11144
rect 12032 11092 12038 11144
rect 12084 11141 12112 11172
rect 12069 11135 12127 11141
rect 12069 11101 12081 11135
rect 12115 11101 12127 11135
rect 12069 11095 12127 11101
rect 12253 11135 12311 11141
rect 12253 11101 12265 11135
rect 12299 11132 12311 11135
rect 12342 11132 12348 11144
rect 12299 11104 12348 11132
rect 12299 11101 12311 11104
rect 12253 11095 12311 11101
rect 12342 11092 12348 11104
rect 12400 11092 12406 11144
rect 12710 11092 12716 11144
rect 12768 11132 12774 11144
rect 12897 11135 12955 11141
rect 12897 11132 12909 11135
rect 12768 11104 12909 11132
rect 12768 11092 12774 11104
rect 12897 11101 12909 11104
rect 12943 11101 12955 11135
rect 13004 11132 13032 11172
rect 13078 11160 13084 11212
rect 13136 11160 13142 11212
rect 13630 11160 13636 11212
rect 13688 11160 13694 11212
rect 15194 11160 15200 11212
rect 15252 11200 15258 11212
rect 16040 11200 16068 11308
rect 16390 11296 16396 11308
rect 16448 11336 16454 11348
rect 17218 11336 17224 11348
rect 16448 11308 17224 11336
rect 16448 11296 16454 11308
rect 17218 11296 17224 11308
rect 17276 11296 17282 11348
rect 18690 11296 18696 11348
rect 18748 11296 18754 11348
rect 19794 11296 19800 11348
rect 19852 11296 19858 11348
rect 19978 11296 19984 11348
rect 20036 11336 20042 11348
rect 21174 11336 21180 11348
rect 20036 11308 21180 11336
rect 20036 11296 20042 11308
rect 21174 11296 21180 11308
rect 21232 11296 21238 11348
rect 21358 11296 21364 11348
rect 21416 11336 21422 11348
rect 21542 11336 21548 11348
rect 21416 11308 21548 11336
rect 21416 11296 21422 11308
rect 21542 11296 21548 11308
rect 21600 11296 21606 11348
rect 23477 11339 23535 11345
rect 23477 11305 23489 11339
rect 23523 11336 23535 11339
rect 24213 11339 24271 11345
rect 23523 11308 23796 11336
rect 23523 11305 23535 11308
rect 23477 11299 23535 11305
rect 17678 11228 17684 11280
rect 17736 11268 17742 11280
rect 18708 11268 18736 11296
rect 20162 11268 20168 11280
rect 17736 11240 20168 11268
rect 17736 11228 17742 11240
rect 20162 11228 20168 11240
rect 20220 11228 20226 11280
rect 21100 11240 23520 11268
rect 15252 11172 15792 11200
rect 15252 11160 15258 11172
rect 15764 11144 15792 11172
rect 15948 11172 16068 11200
rect 16577 11203 16635 11209
rect 13262 11132 13268 11144
rect 13004 11104 13268 11132
rect 12897 11095 12955 11101
rect 13262 11092 13268 11104
rect 13320 11092 13326 11144
rect 13538 11092 13544 11144
rect 13596 11092 13602 11144
rect 13722 11092 13728 11144
rect 13780 11092 13786 11144
rect 15378 11092 15384 11144
rect 15436 11092 15442 11144
rect 15565 11135 15623 11141
rect 15565 11101 15577 11135
rect 15611 11101 15623 11135
rect 15565 11095 15623 11101
rect 2004 11036 4108 11064
rect 2004 11024 2010 11036
rect 4080 10996 4108 11036
rect 5810 11024 5816 11076
rect 5868 11064 5874 11076
rect 6917 11067 6975 11073
rect 6917 11064 6929 11067
rect 5868 11036 6929 11064
rect 5868 11024 5874 11036
rect 6917 11033 6929 11036
rect 6963 11033 6975 11067
rect 9861 11067 9919 11073
rect 6917 11027 6975 11033
rect 8588 11036 9720 11064
rect 4706 10996 4712 11008
rect 4080 10968 4712 10996
rect 4706 10956 4712 10968
rect 4764 10956 4770 11008
rect 5353 10999 5411 11005
rect 5353 10965 5365 10999
rect 5399 10996 5411 10999
rect 6454 10996 6460 11008
rect 5399 10968 6460 10996
rect 5399 10965 5411 10968
rect 5353 10959 5411 10965
rect 6454 10956 6460 10968
rect 6512 10956 6518 11008
rect 6730 10956 6736 11008
rect 6788 10996 6794 11008
rect 8588 10996 8616 11036
rect 6788 10968 8616 10996
rect 6788 10956 6794 10968
rect 8662 10956 8668 11008
rect 8720 10996 8726 11008
rect 9585 10999 9643 11005
rect 9585 10996 9597 10999
rect 8720 10968 9597 10996
rect 8720 10956 8726 10968
rect 9585 10965 9597 10968
rect 9631 10965 9643 10999
rect 9692 10996 9720 11036
rect 9861 11033 9873 11067
rect 9907 11064 9919 11067
rect 10505 11067 10563 11073
rect 10505 11064 10517 11067
rect 9907 11036 10517 11064
rect 9907 11033 9919 11036
rect 9861 11027 9919 11033
rect 10505 11033 10517 11036
rect 10551 11033 10563 11067
rect 10505 11027 10563 11033
rect 10686 11024 10692 11076
rect 10744 11024 10750 11076
rect 10870 11024 10876 11076
rect 10928 11024 10934 11076
rect 11885 11067 11943 11073
rect 11885 11033 11897 11067
rect 11931 11064 11943 11067
rect 13173 11067 13231 11073
rect 13173 11064 13185 11067
rect 11931 11036 13185 11064
rect 11931 11033 11943 11036
rect 11885 11027 11943 11033
rect 13173 11033 13185 11036
rect 13219 11033 13231 11067
rect 13173 11027 13231 11033
rect 13633 11067 13691 11073
rect 13633 11033 13645 11067
rect 13679 11064 13691 11067
rect 13998 11064 14004 11076
rect 13679 11036 14004 11064
rect 13679 11033 13691 11036
rect 13633 11027 13691 11033
rect 13998 11024 14004 11036
rect 14056 11024 14062 11076
rect 15580 11064 15608 11095
rect 15654 11092 15660 11144
rect 15712 11092 15718 11144
rect 15746 11092 15752 11144
rect 15804 11132 15810 11144
rect 15948 11141 15976 11172
rect 16577 11169 16589 11203
rect 16623 11200 16635 11203
rect 16942 11200 16948 11212
rect 16623 11172 16948 11200
rect 16623 11169 16635 11172
rect 16577 11163 16635 11169
rect 16942 11160 16948 11172
rect 17000 11160 17006 11212
rect 15841 11135 15899 11141
rect 15841 11132 15853 11135
rect 15804 11104 15853 11132
rect 15804 11092 15810 11104
rect 15841 11101 15853 11104
rect 15887 11101 15899 11135
rect 15841 11095 15899 11101
rect 15933 11135 15991 11141
rect 15933 11101 15945 11135
rect 15979 11101 15991 11135
rect 15933 11095 15991 11101
rect 16022 11092 16028 11144
rect 16080 11092 16086 11144
rect 16206 11092 16212 11144
rect 16264 11092 16270 11144
rect 16301 11135 16359 11141
rect 16301 11101 16313 11135
rect 16347 11101 16359 11135
rect 17696 11118 17724 11228
rect 18693 11203 18751 11209
rect 18693 11169 18705 11203
rect 18739 11200 18751 11203
rect 19521 11203 19579 11209
rect 19521 11200 19533 11203
rect 18739 11172 19533 11200
rect 18739 11169 18751 11172
rect 18693 11163 18751 11169
rect 19521 11169 19533 11172
rect 19567 11169 19579 11203
rect 19521 11163 19579 11169
rect 16301 11095 16359 11101
rect 16224 11064 16252 11092
rect 15580 11036 16252 11064
rect 16316 11064 16344 11095
rect 18322 11092 18328 11144
rect 18380 11092 18386 11144
rect 19334 11092 19340 11144
rect 19392 11092 19398 11144
rect 19426 11092 19432 11144
rect 19484 11092 19490 11144
rect 19613 11135 19671 11141
rect 19613 11101 19625 11135
rect 19659 11101 19671 11135
rect 19613 11095 19671 11101
rect 16482 11064 16488 11076
rect 16316 11036 16488 11064
rect 16482 11024 16488 11036
rect 16540 11024 16546 11076
rect 18506 11024 18512 11076
rect 18564 11024 18570 11076
rect 18966 11024 18972 11076
rect 19024 11064 19030 11076
rect 19628 11064 19656 11095
rect 19794 11092 19800 11144
rect 19852 11132 19858 11144
rect 20438 11132 20444 11144
rect 19852 11104 20444 11132
rect 19852 11092 19858 11104
rect 20438 11092 20444 11104
rect 20496 11132 20502 11144
rect 21100 11141 21128 11240
rect 21542 11200 21548 11212
rect 21284 11172 21548 11200
rect 21284 11144 21312 11172
rect 21542 11160 21548 11172
rect 21600 11160 21606 11212
rect 21085 11135 21143 11141
rect 21085 11132 21097 11135
rect 20496 11104 21097 11132
rect 20496 11092 20502 11104
rect 21085 11101 21097 11104
rect 21131 11101 21143 11135
rect 21085 11095 21143 11101
rect 21266 11092 21272 11144
rect 21324 11092 21330 11144
rect 21358 11092 21364 11144
rect 21416 11092 21422 11144
rect 21637 11135 21695 11141
rect 21637 11101 21649 11135
rect 21683 11101 21695 11135
rect 21637 11095 21695 11101
rect 19024 11036 19656 11064
rect 19024 11024 19030 11036
rect 20806 11024 20812 11076
rect 20864 11064 20870 11076
rect 21652 11064 21680 11095
rect 23198 11092 23204 11144
rect 23256 11092 23262 11144
rect 23492 11073 23520 11240
rect 23569 11135 23627 11141
rect 23569 11101 23581 11135
rect 23615 11132 23627 11135
rect 23658 11132 23664 11144
rect 23615 11104 23664 11132
rect 23615 11101 23627 11104
rect 23569 11095 23627 11101
rect 23658 11092 23664 11104
rect 23716 11092 23722 11144
rect 23768 11141 23796 11308
rect 24213 11305 24225 11339
rect 24259 11336 24271 11339
rect 24486 11336 24492 11348
rect 24259 11308 24492 11336
rect 24259 11305 24271 11308
rect 24213 11299 24271 11305
rect 24486 11296 24492 11308
rect 24544 11336 24550 11348
rect 24654 11339 24712 11345
rect 24654 11336 24666 11339
rect 24544 11308 24666 11336
rect 24544 11296 24550 11308
rect 24654 11305 24666 11308
rect 24700 11305 24712 11339
rect 24654 11299 24712 11305
rect 24854 11296 24860 11348
rect 24912 11336 24918 11348
rect 26145 11339 26203 11345
rect 26145 11336 26157 11339
rect 24912 11308 26157 11336
rect 24912 11296 24918 11308
rect 26145 11305 26157 11308
rect 26191 11305 26203 11339
rect 26145 11299 26203 11305
rect 23845 11271 23903 11277
rect 23845 11237 23857 11271
rect 23891 11268 23903 11271
rect 23934 11268 23940 11280
rect 23891 11240 23940 11268
rect 23891 11237 23903 11240
rect 23845 11231 23903 11237
rect 23934 11228 23940 11240
rect 23992 11228 23998 11280
rect 24397 11203 24455 11209
rect 24397 11169 24409 11203
rect 24443 11200 24455 11203
rect 24670 11200 24676 11212
rect 24443 11172 24676 11200
rect 24443 11169 24455 11172
rect 24397 11163 24455 11169
rect 24670 11160 24676 11172
rect 24728 11160 24734 11212
rect 23753 11135 23811 11141
rect 23753 11101 23765 11135
rect 23799 11101 23811 11135
rect 23753 11095 23811 11101
rect 23934 11092 23940 11144
rect 23992 11092 23998 11144
rect 24029 11135 24087 11141
rect 24029 11101 24041 11135
rect 24075 11132 24087 11135
rect 24075 11104 24440 11132
rect 24075 11101 24087 11104
rect 24029 11095 24087 11101
rect 20864 11036 21680 11064
rect 23293 11067 23351 11073
rect 20864 11024 20870 11036
rect 23293 11033 23305 11067
rect 23339 11064 23351 11067
rect 23477 11067 23535 11073
rect 23339 11036 23428 11064
rect 23339 11033 23351 11036
rect 23293 11027 23351 11033
rect 11974 10996 11980 11008
rect 9692 10968 11980 10996
rect 9585 10959 9643 10965
rect 11974 10956 11980 10968
rect 12032 10996 12038 11008
rect 12342 10996 12348 11008
rect 12032 10968 12348 10996
rect 12032 10956 12038 10968
rect 12342 10956 12348 10968
rect 12400 10956 12406 11008
rect 12437 10999 12495 11005
rect 12437 10965 12449 10999
rect 12483 10996 12495 10999
rect 12618 10996 12624 11008
rect 12483 10968 12624 10996
rect 12483 10965 12495 10968
rect 12437 10959 12495 10965
rect 12618 10956 12624 10968
rect 12676 10956 12682 11008
rect 12986 10956 12992 11008
rect 13044 10996 13050 11008
rect 13357 10999 13415 11005
rect 13357 10996 13369 10999
rect 13044 10968 13369 10996
rect 13044 10956 13050 10968
rect 13357 10965 13369 10968
rect 13403 10965 13415 10999
rect 13357 10959 13415 10965
rect 16114 10956 16120 11008
rect 16172 10996 16178 11008
rect 16209 10999 16267 11005
rect 16209 10996 16221 10999
rect 16172 10968 16221 10996
rect 16172 10956 16178 10968
rect 16209 10965 16221 10968
rect 16255 10965 16267 10999
rect 16209 10959 16267 10965
rect 16574 10956 16580 11008
rect 16632 10996 16638 11008
rect 17586 10996 17592 11008
rect 16632 10968 17592 10996
rect 16632 10956 16638 10968
rect 17586 10956 17592 10968
rect 17644 10996 17650 11008
rect 18049 10999 18107 11005
rect 18049 10996 18061 10999
rect 17644 10968 18061 10996
rect 17644 10956 17650 10968
rect 18049 10965 18061 10968
rect 18095 10965 18107 10999
rect 18049 10959 18107 10965
rect 20714 10956 20720 11008
rect 20772 10996 20778 11008
rect 20901 10999 20959 11005
rect 20901 10996 20913 10999
rect 20772 10968 20913 10996
rect 20772 10956 20778 10968
rect 20901 10965 20913 10968
rect 20947 10965 20959 10999
rect 23400 10996 23428 11036
rect 23477 11033 23489 11067
rect 23523 11064 23535 11067
rect 24210 11064 24216 11076
rect 23523 11036 24216 11064
rect 23523 11033 23535 11036
rect 23477 11027 23535 11033
rect 24210 11024 24216 11036
rect 24268 11024 24274 11076
rect 24412 11064 24440 11104
rect 24762 11064 24768 11076
rect 24412 11036 24768 11064
rect 24762 11024 24768 11036
rect 24820 11024 24826 11076
rect 25130 11024 25136 11076
rect 25188 11024 25194 11076
rect 24026 10996 24032 11008
rect 23400 10968 24032 10996
rect 20901 10959 20959 10965
rect 24026 10956 24032 10968
rect 24084 10956 24090 11008
rect 1104 10906 28152 10928
rect 1104 10854 4874 10906
rect 4926 10854 4938 10906
rect 4990 10854 5002 10906
rect 5054 10854 5066 10906
rect 5118 10854 5130 10906
rect 5182 10854 28152 10906
rect 1104 10832 28152 10854
rect 3142 10792 3148 10804
rect 2746 10764 3148 10792
rect 2746 10724 2774 10764
rect 3142 10752 3148 10764
rect 3200 10792 3206 10804
rect 3237 10795 3295 10801
rect 3237 10792 3249 10795
rect 3200 10764 3249 10792
rect 3200 10752 3206 10764
rect 3237 10761 3249 10764
rect 3283 10761 3295 10795
rect 3237 10755 3295 10761
rect 5810 10752 5816 10804
rect 5868 10752 5874 10804
rect 8662 10752 8668 10804
rect 8720 10752 8726 10804
rect 9858 10752 9864 10804
rect 9916 10792 9922 10804
rect 9916 10764 13216 10792
rect 9916 10752 9922 10764
rect 6454 10724 6460 10736
rect 2700 10696 2774 10724
rect 6042 10696 6460 10724
rect 1854 10616 1860 10668
rect 1912 10616 1918 10668
rect 2700 10665 2728 10696
rect 2685 10659 2743 10665
rect 2685 10625 2697 10659
rect 2731 10625 2743 10659
rect 2685 10619 2743 10625
rect 3145 10659 3203 10665
rect 3145 10625 3157 10659
rect 3191 10625 3203 10659
rect 3145 10619 3203 10625
rect 3329 10659 3387 10665
rect 3329 10625 3341 10659
rect 3375 10656 3387 10659
rect 3418 10656 3424 10668
rect 3375 10628 3424 10656
rect 3375 10625 3387 10628
rect 3329 10619 3387 10625
rect 1946 10548 1952 10600
rect 2004 10548 2010 10600
rect 2593 10591 2651 10597
rect 2593 10557 2605 10591
rect 2639 10588 2651 10591
rect 2866 10588 2872 10600
rect 2639 10560 2872 10588
rect 2639 10557 2651 10560
rect 2593 10551 2651 10557
rect 2866 10548 2872 10560
rect 2924 10548 2930 10600
rect 2225 10523 2283 10529
rect 2225 10489 2237 10523
rect 2271 10520 2283 10523
rect 2682 10520 2688 10532
rect 2271 10492 2688 10520
rect 2271 10489 2283 10492
rect 2225 10483 2283 10489
rect 2682 10480 2688 10492
rect 2740 10520 2746 10532
rect 3160 10520 3188 10619
rect 3418 10616 3424 10628
rect 3476 10616 3482 10668
rect 6042 10665 6070 10696
rect 6454 10684 6460 10696
rect 6512 10684 6518 10736
rect 8478 10684 8484 10736
rect 8536 10724 8542 10736
rect 9677 10727 9735 10733
rect 8536 10696 8800 10724
rect 8536 10684 8542 10696
rect 6027 10659 6085 10665
rect 6027 10625 6039 10659
rect 6073 10625 6085 10659
rect 6027 10619 6085 10625
rect 6192 10659 6250 10665
rect 6192 10625 6204 10659
rect 6238 10654 6250 10659
rect 6362 10656 6368 10668
rect 6288 10654 6368 10656
rect 6238 10628 6368 10654
rect 6238 10626 6316 10628
rect 6238 10625 6250 10626
rect 6192 10619 6250 10625
rect 6362 10616 6368 10628
rect 6420 10656 6426 10668
rect 6549 10659 6607 10665
rect 6549 10656 6561 10659
rect 6420 10628 6561 10656
rect 6420 10616 6426 10628
rect 6549 10625 6561 10628
rect 6595 10625 6607 10659
rect 6549 10619 6607 10625
rect 7377 10659 7435 10665
rect 7377 10625 7389 10659
rect 7423 10656 7435 10659
rect 8570 10656 8576 10668
rect 7423 10628 8576 10656
rect 7423 10625 7435 10628
rect 7377 10619 7435 10625
rect 8570 10616 8576 10628
rect 8628 10616 8634 10668
rect 8772 10665 8800 10696
rect 9677 10693 9689 10727
rect 9723 10724 9735 10727
rect 9766 10724 9772 10736
rect 9723 10696 9772 10724
rect 9723 10693 9735 10696
rect 9677 10687 9735 10693
rect 9766 10684 9772 10696
rect 9824 10724 9830 10736
rect 10045 10727 10103 10733
rect 10045 10724 10057 10727
rect 9824 10696 10057 10724
rect 9824 10684 9830 10696
rect 10045 10693 10057 10696
rect 10091 10693 10103 10727
rect 10045 10687 10103 10693
rect 11609 10727 11667 10733
rect 11609 10693 11621 10727
rect 11655 10724 11667 10727
rect 11655 10696 11836 10724
rect 11655 10693 11667 10696
rect 11609 10687 11667 10693
rect 11808 10668 11836 10696
rect 8757 10659 8815 10665
rect 8757 10625 8769 10659
rect 8803 10625 8815 10659
rect 8757 10619 8815 10625
rect 9214 10616 9220 10668
rect 9272 10616 9278 10668
rect 9401 10659 9459 10665
rect 9401 10625 9413 10659
rect 9447 10656 9459 10659
rect 9493 10659 9551 10665
rect 9493 10656 9505 10659
rect 9447 10628 9505 10656
rect 9447 10625 9459 10628
rect 9401 10619 9459 10625
rect 9493 10625 9505 10628
rect 9539 10625 9551 10659
rect 9493 10619 9551 10625
rect 9858 10616 9864 10668
rect 9916 10616 9922 10668
rect 9953 10659 10011 10665
rect 9953 10625 9965 10659
rect 9999 10625 10011 10659
rect 9953 10619 10011 10625
rect 10137 10659 10195 10665
rect 10137 10625 10149 10659
rect 10183 10625 10195 10659
rect 10137 10619 10195 10625
rect 6454 10548 6460 10600
rect 6512 10548 6518 10600
rect 7469 10591 7527 10597
rect 7469 10588 7481 10591
rect 6932 10560 7481 10588
rect 6932 10529 6960 10560
rect 7469 10557 7481 10560
rect 7515 10588 7527 10591
rect 7558 10588 7564 10600
rect 7515 10560 7564 10588
rect 7515 10557 7527 10560
rect 7469 10551 7527 10557
rect 7558 10548 7564 10560
rect 7616 10548 7622 10600
rect 8386 10548 8392 10600
rect 8444 10588 8450 10600
rect 9033 10591 9091 10597
rect 9033 10588 9045 10591
rect 8444 10560 9045 10588
rect 8444 10548 8450 10560
rect 9033 10557 9045 10560
rect 9079 10557 9091 10591
rect 9232 10588 9260 10616
rect 9968 10588 9996 10619
rect 9232 10560 9996 10588
rect 9033 10551 9091 10557
rect 2740 10492 3188 10520
rect 6917 10523 6975 10529
rect 2740 10480 2746 10492
rect 6917 10489 6929 10523
rect 6963 10489 6975 10523
rect 6917 10483 6975 10489
rect 7745 10523 7803 10529
rect 7745 10489 7757 10523
rect 7791 10520 7803 10523
rect 8846 10520 8852 10532
rect 7791 10492 8852 10520
rect 7791 10489 7803 10492
rect 7745 10483 7803 10489
rect 8846 10480 8852 10492
rect 8904 10480 8910 10532
rect 9048 10520 9076 10551
rect 10152 10520 10180 10619
rect 10410 10616 10416 10668
rect 10468 10656 10474 10668
rect 11514 10656 11520 10668
rect 10468 10628 11520 10656
rect 10468 10616 10474 10628
rect 11514 10616 11520 10628
rect 11572 10616 11578 10668
rect 11701 10659 11759 10665
rect 11701 10625 11713 10659
rect 11747 10625 11759 10659
rect 11701 10619 11759 10625
rect 11422 10548 11428 10600
rect 11480 10588 11486 10600
rect 11716 10588 11744 10619
rect 11790 10616 11796 10668
rect 11848 10616 11854 10668
rect 11882 10616 11888 10668
rect 11940 10616 11946 10668
rect 11974 10616 11980 10668
rect 12032 10656 12038 10668
rect 12069 10659 12127 10665
rect 12069 10656 12081 10659
rect 12032 10628 12081 10656
rect 12032 10616 12038 10628
rect 12069 10625 12081 10628
rect 12115 10625 12127 10659
rect 12069 10619 12127 10625
rect 12158 10616 12164 10668
rect 12216 10616 12222 10668
rect 12345 10659 12403 10665
rect 12345 10625 12357 10659
rect 12391 10656 12403 10659
rect 12391 10628 12572 10656
rect 12391 10625 12403 10628
rect 12345 10619 12403 10625
rect 11480 10560 11744 10588
rect 12544 10588 12572 10628
rect 12618 10616 12624 10668
rect 12676 10616 12682 10668
rect 12802 10616 12808 10668
rect 12860 10616 12866 10668
rect 12986 10616 12992 10668
rect 13044 10616 13050 10668
rect 13188 10665 13216 10764
rect 15470 10752 15476 10804
rect 15528 10752 15534 10804
rect 16298 10752 16304 10804
rect 16356 10792 16362 10804
rect 16393 10795 16451 10801
rect 16393 10792 16405 10795
rect 16356 10764 16405 10792
rect 16356 10752 16362 10764
rect 16393 10761 16405 10764
rect 16439 10761 16451 10795
rect 16393 10755 16451 10761
rect 18138 10752 18144 10804
rect 18196 10752 18202 10804
rect 18414 10752 18420 10804
rect 18472 10792 18478 10804
rect 18782 10792 18788 10804
rect 18472 10764 18788 10792
rect 18472 10752 18478 10764
rect 18782 10752 18788 10764
rect 18840 10792 18846 10804
rect 18840 10764 21220 10792
rect 18840 10752 18846 10764
rect 15930 10684 15936 10736
rect 15988 10724 15994 10736
rect 16025 10727 16083 10733
rect 16025 10724 16037 10727
rect 15988 10696 16037 10724
rect 15988 10684 15994 10696
rect 16025 10693 16037 10696
rect 16071 10693 16083 10727
rect 17405 10727 17463 10733
rect 16025 10687 16083 10693
rect 16132 10696 16988 10724
rect 16132 10668 16160 10696
rect 13173 10659 13231 10665
rect 13173 10625 13185 10659
rect 13219 10625 13231 10659
rect 13173 10619 13231 10625
rect 13998 10616 14004 10668
rect 14056 10616 14062 10668
rect 14185 10659 14243 10665
rect 14185 10625 14197 10659
rect 14231 10625 14243 10659
rect 14185 10619 14243 10625
rect 12897 10591 12955 10597
rect 12897 10588 12909 10591
rect 12544 10560 12909 10588
rect 11480 10548 11486 10560
rect 12897 10557 12909 10560
rect 12943 10588 12955 10591
rect 13262 10588 13268 10600
rect 12943 10560 13268 10588
rect 12943 10557 12955 10560
rect 12897 10551 12955 10557
rect 13262 10548 13268 10560
rect 13320 10548 13326 10600
rect 13357 10591 13415 10597
rect 13357 10557 13369 10591
rect 13403 10588 13415 10591
rect 14200 10588 14228 10619
rect 14458 10616 14464 10668
rect 14516 10616 14522 10668
rect 14734 10616 14740 10668
rect 14792 10656 14798 10668
rect 15105 10659 15163 10665
rect 15105 10656 15117 10659
rect 14792 10628 15117 10656
rect 14792 10616 14798 10628
rect 15105 10625 15117 10628
rect 15151 10625 15163 10659
rect 15105 10619 15163 10625
rect 15289 10659 15347 10665
rect 15289 10625 15301 10659
rect 15335 10656 15347 10659
rect 16114 10656 16120 10668
rect 15335 10628 16120 10656
rect 15335 10625 15347 10628
rect 15289 10619 15347 10625
rect 16114 10616 16120 10628
rect 16172 10616 16178 10668
rect 16209 10659 16267 10665
rect 16209 10625 16221 10659
rect 16255 10625 16267 10659
rect 16209 10619 16267 10625
rect 15470 10588 15476 10600
rect 13403 10560 14228 10588
rect 14292 10560 15476 10588
rect 13403 10557 13415 10560
rect 13357 10551 13415 10557
rect 9048 10492 10180 10520
rect 10686 10480 10692 10532
rect 10744 10520 10750 10532
rect 14090 10520 14096 10532
rect 10744 10492 14096 10520
rect 10744 10480 10750 10492
rect 14090 10480 14096 10492
rect 14148 10480 14154 10532
rect 3053 10455 3111 10461
rect 3053 10421 3065 10455
rect 3099 10452 3111 10455
rect 4062 10452 4068 10464
rect 3099 10424 4068 10452
rect 3099 10421 3111 10424
rect 3053 10415 3111 10421
rect 4062 10412 4068 10424
rect 4120 10412 4126 10464
rect 5350 10412 5356 10464
rect 5408 10452 5414 10464
rect 10410 10452 10416 10464
rect 5408 10424 10416 10452
rect 5408 10412 5414 10424
rect 10410 10412 10416 10424
rect 10468 10412 10474 10464
rect 12618 10412 12624 10464
rect 12676 10452 12682 10464
rect 13446 10452 13452 10464
rect 12676 10424 13452 10452
rect 12676 10412 12682 10424
rect 13446 10412 13452 10424
rect 13504 10452 13510 10464
rect 14292 10452 14320 10560
rect 15470 10548 15476 10560
rect 15528 10588 15534 10600
rect 16224 10588 16252 10619
rect 16298 10616 16304 10668
rect 16356 10656 16362 10668
rect 16485 10659 16543 10665
rect 16485 10658 16497 10659
rect 16408 10656 16497 10658
rect 16356 10630 16497 10656
rect 16356 10628 16436 10630
rect 16356 10616 16362 10628
rect 16485 10625 16497 10630
rect 16531 10625 16543 10659
rect 16485 10619 16543 10625
rect 16666 10616 16672 10668
rect 16724 10616 16730 10668
rect 16853 10659 16911 10665
rect 16853 10625 16865 10659
rect 16899 10658 16911 10659
rect 16960 10658 16988 10696
rect 17405 10693 17417 10727
rect 17451 10724 17463 10727
rect 18506 10724 18512 10736
rect 17451 10696 18512 10724
rect 17451 10693 17463 10696
rect 17405 10687 17463 10693
rect 18506 10684 18512 10696
rect 18564 10684 18570 10736
rect 20809 10727 20867 10733
rect 20809 10693 20821 10727
rect 20855 10724 20867 10727
rect 20993 10727 21051 10733
rect 20993 10724 21005 10727
rect 20855 10696 21005 10724
rect 20855 10693 20867 10696
rect 20809 10687 20867 10693
rect 20993 10693 21005 10696
rect 21039 10693 21051 10727
rect 21192 10724 21220 10764
rect 23842 10752 23848 10804
rect 23900 10792 23906 10804
rect 24486 10792 24492 10804
rect 24544 10801 24550 10804
rect 24544 10795 24563 10801
rect 23900 10764 24492 10792
rect 23900 10752 23906 10764
rect 24486 10752 24492 10764
rect 24551 10761 24563 10795
rect 24544 10755 24563 10761
rect 24544 10752 24550 10755
rect 21726 10724 21732 10736
rect 21192 10696 21312 10724
rect 20993 10687 21051 10693
rect 16899 10630 16988 10658
rect 16899 10625 16911 10630
rect 16853 10619 16911 10625
rect 17218 10616 17224 10668
rect 17276 10616 17282 10668
rect 17494 10616 17500 10668
rect 17552 10616 17558 10668
rect 17586 10616 17592 10668
rect 17644 10656 17650 10668
rect 17644 10628 17689 10656
rect 17644 10616 17650 10628
rect 17770 10616 17776 10668
rect 17828 10616 17834 10668
rect 17862 10616 17868 10668
rect 17920 10616 17926 10668
rect 17962 10659 18020 10665
rect 17962 10625 17974 10659
rect 18008 10656 18020 10659
rect 18138 10656 18144 10668
rect 18008 10628 18144 10656
rect 18008 10625 18020 10628
rect 17962 10619 18020 10625
rect 18138 10616 18144 10628
rect 18196 10616 18202 10668
rect 19886 10616 19892 10668
rect 19944 10656 19950 10668
rect 20165 10659 20223 10665
rect 20165 10656 20177 10659
rect 19944 10628 20177 10656
rect 19944 10616 19950 10628
rect 20165 10625 20177 10628
rect 20211 10656 20223 10659
rect 20441 10659 20499 10665
rect 20441 10656 20453 10659
rect 20211 10628 20453 10656
rect 20211 10625 20223 10628
rect 20165 10619 20223 10625
rect 20441 10625 20453 10628
rect 20487 10625 20499 10659
rect 20441 10619 20499 10625
rect 20625 10659 20683 10665
rect 20625 10625 20637 10659
rect 20671 10656 20683 10659
rect 20714 10656 20720 10668
rect 20671 10628 20720 10656
rect 20671 10625 20683 10628
rect 20625 10619 20683 10625
rect 20714 10616 20720 10628
rect 20772 10616 20778 10668
rect 20901 10659 20959 10665
rect 20901 10625 20913 10659
rect 20947 10625 20959 10659
rect 20901 10619 20959 10625
rect 15528 10560 16252 10588
rect 16939 10591 16997 10597
rect 15528 10548 15534 10560
rect 16939 10557 16951 10591
rect 16985 10557 16997 10591
rect 16939 10551 16997 10557
rect 17037 10591 17095 10597
rect 17037 10557 17049 10591
rect 17083 10557 17095 10591
rect 20916 10588 20944 10619
rect 21174 10616 21180 10668
rect 21232 10616 21238 10668
rect 21284 10665 21312 10696
rect 21468 10696 21732 10724
rect 21468 10665 21496 10696
rect 21726 10684 21732 10696
rect 21784 10684 21790 10736
rect 23750 10684 23756 10736
rect 23808 10684 23814 10736
rect 24118 10684 24124 10736
rect 24176 10724 24182 10736
rect 24305 10727 24363 10733
rect 24305 10724 24317 10727
rect 24176 10696 24317 10724
rect 24176 10684 24182 10696
rect 24305 10693 24317 10696
rect 24351 10693 24363 10727
rect 24305 10687 24363 10693
rect 24394 10684 24400 10736
rect 24452 10724 24458 10736
rect 25133 10727 25191 10733
rect 25133 10724 25145 10727
rect 24452 10696 25145 10724
rect 24452 10684 24458 10696
rect 25133 10693 25145 10696
rect 25179 10693 25191 10727
rect 25133 10687 25191 10693
rect 21269 10659 21327 10665
rect 21269 10625 21281 10659
rect 21315 10625 21327 10659
rect 21269 10619 21327 10625
rect 21453 10659 21511 10665
rect 21453 10625 21465 10659
rect 21499 10625 21511 10659
rect 21453 10619 21511 10625
rect 21542 10616 21548 10668
rect 21600 10616 21606 10668
rect 24026 10616 24032 10668
rect 24084 10616 24090 10668
rect 24578 10656 24584 10668
rect 24228 10628 24584 10656
rect 21818 10588 21824 10600
rect 20916 10560 21824 10588
rect 17037 10551 17095 10557
rect 14645 10523 14703 10529
rect 14645 10489 14657 10523
rect 14691 10520 14703 10523
rect 16960 10520 16988 10551
rect 14691 10492 16988 10520
rect 14691 10489 14703 10492
rect 14645 10483 14703 10489
rect 13504 10424 14320 10452
rect 13504 10412 13510 10424
rect 14458 10412 14464 10464
rect 14516 10452 14522 10464
rect 15105 10455 15163 10461
rect 15105 10452 15117 10455
rect 14516 10424 15117 10452
rect 14516 10412 14522 10424
rect 15105 10421 15117 10424
rect 15151 10421 15163 10455
rect 15105 10415 15163 10421
rect 16022 10412 16028 10464
rect 16080 10452 16086 10464
rect 16390 10452 16396 10464
rect 16080 10424 16396 10452
rect 16080 10412 16086 10424
rect 16390 10412 16396 10424
rect 16448 10452 16454 10464
rect 17052 10452 17080 10551
rect 21818 10548 21824 10560
rect 21876 10548 21882 10600
rect 21910 10548 21916 10600
rect 21968 10588 21974 10600
rect 23845 10591 23903 10597
rect 23845 10588 23857 10591
rect 21968 10560 23857 10588
rect 21968 10548 21974 10560
rect 23845 10557 23857 10560
rect 23891 10557 23903 10591
rect 23845 10551 23903 10557
rect 18598 10480 18604 10532
rect 18656 10520 18662 10532
rect 20898 10520 20904 10532
rect 18656 10492 20904 10520
rect 18656 10480 18662 10492
rect 20898 10480 20904 10492
rect 20956 10520 20962 10532
rect 21726 10520 21732 10532
rect 20956 10492 21732 10520
rect 20956 10480 20962 10492
rect 21726 10480 21732 10492
rect 21784 10480 21790 10532
rect 23658 10480 23664 10532
rect 23716 10520 23722 10532
rect 24228 10529 24256 10628
rect 24578 10616 24584 10628
rect 24636 10656 24642 10668
rect 24765 10659 24823 10665
rect 24765 10656 24777 10659
rect 24636 10628 24777 10656
rect 24636 10616 24642 10628
rect 24765 10625 24777 10628
rect 24811 10625 24823 10659
rect 24765 10619 24823 10625
rect 24949 10659 25007 10665
rect 24949 10625 24961 10659
rect 24995 10625 25007 10659
rect 24949 10619 25007 10625
rect 24213 10523 24271 10529
rect 24213 10520 24225 10523
rect 23716 10492 24225 10520
rect 23716 10480 23722 10492
rect 24213 10489 24225 10492
rect 24259 10489 24271 10523
rect 24213 10483 24271 10489
rect 24762 10480 24768 10532
rect 24820 10520 24826 10532
rect 24964 10520 24992 10619
rect 24820 10492 24992 10520
rect 24820 10480 24826 10492
rect 16448 10424 17080 10452
rect 16448 10412 16454 10424
rect 20254 10412 20260 10464
rect 20312 10412 20318 10464
rect 23198 10412 23204 10464
rect 23256 10452 23262 10464
rect 23842 10452 23848 10464
rect 23256 10424 23848 10452
rect 23256 10412 23262 10424
rect 23842 10412 23848 10424
rect 23900 10412 23906 10464
rect 24394 10412 24400 10464
rect 24452 10452 24458 10464
rect 24489 10455 24547 10461
rect 24489 10452 24501 10455
rect 24452 10424 24501 10452
rect 24452 10412 24458 10424
rect 24489 10421 24501 10424
rect 24535 10421 24547 10455
rect 24489 10415 24547 10421
rect 24673 10455 24731 10461
rect 24673 10421 24685 10455
rect 24719 10452 24731 10455
rect 24946 10452 24952 10464
rect 24719 10424 24952 10452
rect 24719 10421 24731 10424
rect 24673 10415 24731 10421
rect 24946 10412 24952 10424
rect 25004 10412 25010 10464
rect 1104 10362 28152 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 28152 10362
rect 1104 10288 28152 10310
rect 7745 10251 7803 10257
rect 7745 10217 7757 10251
rect 7791 10248 7803 10251
rect 8386 10248 8392 10260
rect 7791 10220 8392 10248
rect 7791 10217 7803 10220
rect 7745 10211 7803 10217
rect 8386 10208 8392 10220
rect 8444 10208 8450 10260
rect 8481 10251 8539 10257
rect 8481 10217 8493 10251
rect 8527 10248 8539 10251
rect 8662 10248 8668 10260
rect 8527 10220 8668 10248
rect 8527 10217 8539 10220
rect 8481 10211 8539 10217
rect 3145 10183 3203 10189
rect 3145 10149 3157 10183
rect 3191 10180 3203 10183
rect 4614 10180 4620 10192
rect 3191 10152 4620 10180
rect 3191 10149 3203 10152
rect 3145 10143 3203 10149
rect 4614 10140 4620 10152
rect 4672 10140 4678 10192
rect 8294 10180 8300 10192
rect 7944 10152 8300 10180
rect 2682 10072 2688 10124
rect 2740 10072 2746 10124
rect 4062 10072 4068 10124
rect 4120 10072 4126 10124
rect 5350 10112 5356 10124
rect 4448 10084 5356 10112
rect 2777 10047 2835 10053
rect 2777 10013 2789 10047
rect 2823 10044 2835 10047
rect 3418 10044 3424 10056
rect 2823 10016 3424 10044
rect 2823 10013 2835 10016
rect 2777 10007 2835 10013
rect 3418 10004 3424 10016
rect 3476 10004 3482 10056
rect 4448 10053 4476 10084
rect 5350 10072 5356 10084
rect 5408 10072 5414 10124
rect 5442 10072 5448 10124
rect 5500 10112 5506 10124
rect 7944 10121 7972 10152
rect 8294 10140 8300 10152
rect 8352 10140 8358 10192
rect 7929 10115 7987 10121
rect 8496 10120 8524 10211
rect 8662 10208 8668 10220
rect 8720 10208 8726 10260
rect 11882 10208 11888 10260
rect 11940 10248 11946 10260
rect 12161 10251 12219 10257
rect 12161 10248 12173 10251
rect 11940 10220 12173 10248
rect 11940 10208 11946 10220
rect 12161 10217 12173 10220
rect 12207 10217 12219 10251
rect 12986 10248 12992 10260
rect 12161 10211 12219 10217
rect 12406 10220 12992 10248
rect 12406 10180 12434 10220
rect 12986 10208 12992 10220
rect 13044 10208 13050 10260
rect 13078 10208 13084 10260
rect 13136 10248 13142 10260
rect 13173 10251 13231 10257
rect 13173 10248 13185 10251
rect 13136 10220 13185 10248
rect 13136 10208 13142 10220
rect 13173 10217 13185 10220
rect 13219 10217 13231 10251
rect 13173 10211 13231 10217
rect 13262 10208 13268 10260
rect 13320 10248 13326 10260
rect 14185 10251 14243 10257
rect 14185 10248 14197 10251
rect 13320 10220 14197 10248
rect 13320 10208 13326 10220
rect 14185 10217 14197 10220
rect 14231 10217 14243 10251
rect 14185 10211 14243 10217
rect 14734 10208 14740 10260
rect 14792 10208 14798 10260
rect 16390 10208 16396 10260
rect 16448 10208 16454 10260
rect 16666 10208 16672 10260
rect 16724 10248 16730 10260
rect 16945 10251 17003 10257
rect 16945 10248 16957 10251
rect 16724 10220 16957 10248
rect 16724 10208 16730 10220
rect 16945 10217 16957 10220
rect 16991 10217 17003 10251
rect 16945 10211 17003 10217
rect 20441 10251 20499 10257
rect 20441 10217 20453 10251
rect 20487 10248 20499 10251
rect 22186 10248 22192 10260
rect 20487 10220 22192 10248
rect 20487 10217 20499 10220
rect 20441 10211 20499 10217
rect 22186 10208 22192 10220
rect 22244 10208 22250 10260
rect 24486 10208 24492 10260
rect 24544 10208 24550 10260
rect 24762 10208 24768 10260
rect 24820 10248 24826 10260
rect 24857 10251 24915 10257
rect 24857 10248 24869 10251
rect 24820 10220 24869 10248
rect 24820 10208 24826 10220
rect 24857 10217 24869 10220
rect 24903 10217 24915 10251
rect 24857 10211 24915 10217
rect 11900 10152 12434 10180
rect 13004 10180 13032 10208
rect 13538 10180 13544 10192
rect 13004 10152 13544 10180
rect 7929 10112 7941 10115
rect 5500 10084 7941 10112
rect 5500 10072 5506 10084
rect 7929 10081 7941 10084
rect 7975 10081 7987 10115
rect 8404 10112 8524 10120
rect 7929 10075 7987 10081
rect 8220 10092 8524 10112
rect 8220 10084 8432 10092
rect 3973 10047 4031 10053
rect 3973 10013 3985 10047
rect 4019 10013 4031 10047
rect 3973 10007 4031 10013
rect 4433 10047 4491 10053
rect 4433 10013 4445 10047
rect 4479 10013 4491 10047
rect 4433 10007 4491 10013
rect 4617 10047 4675 10053
rect 4617 10013 4629 10047
rect 4663 10044 4675 10047
rect 4706 10044 4712 10056
rect 4663 10016 4712 10044
rect 4663 10013 4675 10016
rect 4617 10007 4675 10013
rect 3988 9976 4016 10007
rect 4706 10004 4712 10016
rect 4764 10044 4770 10056
rect 5534 10044 5540 10056
rect 4764 10016 5540 10044
rect 4764 10004 4770 10016
rect 5534 10004 5540 10016
rect 5592 10044 5598 10056
rect 6730 10044 6736 10056
rect 5592 10016 6736 10044
rect 5592 10004 5598 10016
rect 6730 10004 6736 10016
rect 6788 10004 6794 10056
rect 8220 10053 8248 10084
rect 8846 10072 8852 10124
rect 8904 10112 8910 10124
rect 8941 10115 8999 10121
rect 8941 10112 8953 10115
rect 8904 10084 8953 10112
rect 8904 10072 8910 10084
rect 8941 10081 8953 10084
rect 8987 10081 8999 10115
rect 8941 10075 8999 10081
rect 7653 10047 7711 10053
rect 7653 10013 7665 10047
rect 7699 10013 7711 10047
rect 7653 10007 7711 10013
rect 7837 10047 7895 10053
rect 7837 10013 7849 10047
rect 7883 10044 7895 10047
rect 8113 10047 8171 10053
rect 7883 10016 8064 10044
rect 7883 10013 7895 10016
rect 7837 10007 7895 10013
rect 4525 9979 4583 9985
rect 4525 9976 4537 9979
rect 3988 9948 4537 9976
rect 4525 9945 4537 9948
rect 4571 9945 4583 9979
rect 7668 9976 7696 10007
rect 7929 9979 7987 9985
rect 7929 9976 7941 9979
rect 7668 9948 7941 9976
rect 4525 9939 4583 9945
rect 7929 9945 7941 9948
rect 7975 9945 7987 9979
rect 7929 9939 7987 9945
rect 4341 9911 4399 9917
rect 4341 9877 4353 9911
rect 4387 9908 4399 9911
rect 4798 9908 4804 9920
rect 4387 9880 4804 9908
rect 4387 9877 4399 9880
rect 4341 9871 4399 9877
rect 4798 9868 4804 9880
rect 4856 9868 4862 9920
rect 8036 9908 8064 10016
rect 8113 10013 8125 10047
rect 8159 10013 8171 10047
rect 8113 10007 8171 10013
rect 8205 10047 8263 10053
rect 8205 10013 8217 10047
rect 8251 10013 8263 10047
rect 8205 10007 8263 10013
rect 8297 10025 8355 10031
rect 8128 9976 8156 10007
rect 8297 9991 8309 10025
rect 8343 9991 8355 10025
rect 8386 10004 8392 10056
rect 8444 10004 8450 10056
rect 9030 10004 9036 10056
rect 9088 10044 9094 10056
rect 9309 10047 9367 10053
rect 9309 10044 9321 10047
rect 9088 10016 9321 10044
rect 9088 10004 9094 10016
rect 9309 10013 9321 10016
rect 9355 10013 9367 10047
rect 9309 10007 9367 10013
rect 9490 10004 9496 10056
rect 9548 10004 9554 10056
rect 9674 10004 9680 10056
rect 9732 10044 9738 10056
rect 9769 10047 9827 10053
rect 9769 10044 9781 10047
rect 9732 10016 9781 10044
rect 9732 10004 9738 10016
rect 9769 10013 9781 10016
rect 9815 10013 9827 10047
rect 9769 10007 9827 10013
rect 11606 10004 11612 10056
rect 11664 10004 11670 10056
rect 11793 10047 11851 10053
rect 11793 10013 11805 10047
rect 11839 10044 11851 10047
rect 11900 10044 11928 10152
rect 13538 10140 13544 10152
rect 13596 10140 13602 10192
rect 14090 10140 14096 10192
rect 14148 10180 14154 10192
rect 16758 10180 16764 10192
rect 14148 10152 15884 10180
rect 14148 10140 14154 10152
rect 12158 10072 12164 10124
rect 12216 10112 12222 10124
rect 13817 10115 13875 10121
rect 13817 10112 13829 10115
rect 12216 10084 13829 10112
rect 12216 10072 12222 10084
rect 13817 10081 13829 10084
rect 13863 10081 13875 10115
rect 13817 10075 13875 10081
rect 13998 10072 14004 10124
rect 14056 10112 14062 10124
rect 14056 10084 14596 10112
rect 14056 10072 14062 10084
rect 11839 10016 11928 10044
rect 11977 10047 12035 10053
rect 11839 10013 11851 10016
rect 11793 10007 11851 10013
rect 11977 10013 11989 10047
rect 12023 10013 12035 10047
rect 11977 10007 12035 10013
rect 8297 9988 8355 9991
rect 8294 9976 8300 9988
rect 8128 9948 8300 9976
rect 8294 9936 8300 9948
rect 8352 9936 8358 9988
rect 9582 9936 9588 9988
rect 9640 9936 9646 9988
rect 8665 9911 8723 9917
rect 8665 9908 8677 9911
rect 8036 9880 8677 9908
rect 8665 9877 8677 9880
rect 8711 9908 8723 9911
rect 8754 9908 8760 9920
rect 8711 9880 8760 9908
rect 8711 9877 8723 9880
rect 8665 9871 8723 9877
rect 8754 9868 8760 9880
rect 8812 9868 8818 9920
rect 9309 9911 9367 9917
rect 9309 9877 9321 9911
rect 9355 9908 9367 9911
rect 9692 9908 9720 10004
rect 9953 9979 10011 9985
rect 9953 9945 9965 9979
rect 9999 9976 10011 9979
rect 11146 9976 11152 9988
rect 9999 9948 11152 9976
rect 9999 9945 10011 9948
rect 9953 9939 10011 9945
rect 11146 9936 11152 9948
rect 11204 9936 11210 9988
rect 11514 9936 11520 9988
rect 11572 9976 11578 9988
rect 11885 9979 11943 9985
rect 11885 9976 11897 9979
rect 11572 9948 11897 9976
rect 11572 9936 11578 9948
rect 11885 9945 11897 9948
rect 11931 9945 11943 9979
rect 11885 9939 11943 9945
rect 11992 9976 12020 10007
rect 12066 10004 12072 10056
rect 12124 10044 12130 10056
rect 12253 10047 12311 10053
rect 12253 10044 12265 10047
rect 12124 10016 12265 10044
rect 12124 10004 12130 10016
rect 12253 10013 12265 10016
rect 12299 10013 12311 10047
rect 12253 10007 12311 10013
rect 12437 10047 12495 10053
rect 12437 10013 12449 10047
rect 12483 10044 12495 10047
rect 12618 10044 12624 10056
rect 12483 10016 12624 10044
rect 12483 10013 12495 10016
rect 12437 10007 12495 10013
rect 12618 10004 12624 10016
rect 12676 10004 12682 10056
rect 12710 10004 12716 10056
rect 12768 10004 12774 10056
rect 12894 10004 12900 10056
rect 12952 10044 12958 10056
rect 13265 10047 13323 10053
rect 13265 10044 13277 10047
rect 12952 10016 13277 10044
rect 12952 10004 12958 10016
rect 13265 10013 13277 10016
rect 13311 10013 13323 10047
rect 13265 10007 13323 10013
rect 13446 10004 13452 10056
rect 13504 10004 13510 10056
rect 13538 10004 13544 10056
rect 13596 10044 13602 10056
rect 13725 10047 13783 10053
rect 13725 10044 13737 10047
rect 13596 10016 13737 10044
rect 13596 10004 13602 10016
rect 13725 10013 13737 10016
rect 13771 10013 13783 10047
rect 13725 10007 13783 10013
rect 14366 10004 14372 10056
rect 14424 10004 14430 10056
rect 14568 10053 14596 10084
rect 14553 10047 14611 10053
rect 14553 10013 14565 10047
rect 14599 10013 14611 10047
rect 15856 10044 15884 10152
rect 16500 10152 16764 10180
rect 16500 10053 16528 10152
rect 16758 10140 16764 10152
rect 16816 10180 16822 10192
rect 17770 10180 17776 10192
rect 16816 10152 17776 10180
rect 16816 10140 16822 10152
rect 17770 10140 17776 10152
rect 17828 10140 17834 10192
rect 18322 10140 18328 10192
rect 18380 10180 18386 10192
rect 18693 10183 18751 10189
rect 18693 10180 18705 10183
rect 18380 10152 18705 10180
rect 18380 10140 18386 10152
rect 18693 10149 18705 10152
rect 18739 10149 18751 10183
rect 18693 10143 18751 10149
rect 19610 10140 19616 10192
rect 19668 10180 19674 10192
rect 24780 10180 24808 10208
rect 19668 10152 19932 10180
rect 19668 10140 19674 10152
rect 16669 10115 16727 10121
rect 16669 10081 16681 10115
rect 16715 10112 16727 10115
rect 17218 10112 17224 10124
rect 16715 10084 17224 10112
rect 16715 10081 16727 10084
rect 16669 10075 16727 10081
rect 17218 10072 17224 10084
rect 17276 10072 17282 10124
rect 17402 10072 17408 10124
rect 17460 10112 17466 10124
rect 18138 10112 18144 10124
rect 17460 10084 18144 10112
rect 17460 10072 17466 10084
rect 18138 10072 18144 10084
rect 18196 10112 18202 10124
rect 18417 10115 18475 10121
rect 18417 10112 18429 10115
rect 18196 10084 18429 10112
rect 18196 10072 18202 10084
rect 18417 10081 18429 10084
rect 18463 10081 18475 10115
rect 18417 10075 18475 10081
rect 18601 10115 18659 10121
rect 18601 10081 18613 10115
rect 18647 10112 18659 10115
rect 19426 10112 19432 10124
rect 18647 10084 19432 10112
rect 18647 10081 18659 10084
rect 18601 10075 18659 10081
rect 19426 10072 19432 10084
rect 19484 10112 19490 10124
rect 19797 10115 19855 10121
rect 19797 10112 19809 10115
rect 19484 10084 19809 10112
rect 19484 10072 19490 10084
rect 19797 10081 19809 10084
rect 19843 10081 19855 10115
rect 19797 10075 19855 10081
rect 16485 10047 16543 10053
rect 16485 10044 16497 10047
rect 15856 10016 16497 10044
rect 14553 10007 14611 10013
rect 16485 10013 16497 10016
rect 16531 10013 16543 10047
rect 16485 10007 16543 10013
rect 16574 10004 16580 10056
rect 16632 10044 16638 10056
rect 16761 10047 16819 10053
rect 16761 10044 16773 10047
rect 16632 10016 16773 10044
rect 16632 10004 16638 10016
rect 16761 10013 16773 10016
rect 16807 10013 16819 10047
rect 16761 10007 16819 10013
rect 16853 10047 16911 10053
rect 16853 10013 16865 10047
rect 16899 10044 16911 10047
rect 16942 10044 16948 10056
rect 16899 10016 16948 10044
rect 16899 10013 16911 10016
rect 16853 10007 16911 10013
rect 16942 10004 16948 10016
rect 17000 10004 17006 10056
rect 17047 10047 17105 10053
rect 17047 10013 17059 10047
rect 17093 10044 17105 10047
rect 17093 10016 17172 10044
rect 17093 10013 17105 10016
rect 17047 10007 17105 10013
rect 12805 9979 12863 9985
rect 12805 9976 12817 9979
rect 11992 9948 12817 9976
rect 9355 9880 9720 9908
rect 9355 9877 9367 9880
rect 9309 9871 9367 9877
rect 11422 9868 11428 9920
rect 11480 9908 11486 9920
rect 11992 9908 12020 9948
rect 12805 9945 12817 9948
rect 12851 9945 12863 9979
rect 12805 9939 12863 9945
rect 13021 9979 13079 9985
rect 13021 9945 13033 9979
rect 13067 9976 13079 9979
rect 13464 9976 13492 10004
rect 13067 9948 13492 9976
rect 13067 9945 13079 9948
rect 13021 9939 13079 9945
rect 14090 9936 14096 9988
rect 14148 9936 14154 9988
rect 15470 9936 15476 9988
rect 15528 9976 15534 9988
rect 17144 9976 17172 10016
rect 18322 10004 18328 10056
rect 18380 10004 18386 10056
rect 18782 10004 18788 10056
rect 18840 10004 18846 10056
rect 19904 10053 19932 10152
rect 24412 10152 24808 10180
rect 20254 10072 20260 10124
rect 20312 10112 20318 10124
rect 20809 10115 20867 10121
rect 20809 10112 20821 10115
rect 20312 10084 20821 10112
rect 20312 10072 20318 10084
rect 20809 10081 20821 10084
rect 20855 10081 20867 10115
rect 20809 10075 20867 10081
rect 19705 10047 19763 10053
rect 19705 10044 19717 10047
rect 19444 10016 19717 10044
rect 17402 9976 17408 9988
rect 15528 9948 16988 9976
rect 17144 9948 17408 9976
rect 15528 9936 15534 9948
rect 11480 9880 12020 9908
rect 11480 9868 11486 9880
rect 12158 9868 12164 9920
rect 12216 9908 12222 9920
rect 12618 9908 12624 9920
rect 12216 9880 12624 9908
rect 12216 9868 12222 9880
rect 12618 9868 12624 9880
rect 12676 9868 12682 9920
rect 12710 9868 12716 9920
rect 12768 9908 12774 9920
rect 13906 9908 13912 9920
rect 12768 9880 13912 9908
rect 12768 9868 12774 9880
rect 13906 9868 13912 9880
rect 13964 9908 13970 9920
rect 16298 9908 16304 9920
rect 13964 9880 16304 9908
rect 13964 9868 13970 9880
rect 16298 9868 16304 9880
rect 16356 9868 16362 9920
rect 16960 9908 16988 9948
rect 17402 9936 17408 9948
rect 17460 9936 17466 9988
rect 18693 9979 18751 9985
rect 18693 9945 18705 9979
rect 18739 9976 18751 9979
rect 19058 9976 19064 9988
rect 18739 9948 19064 9976
rect 18739 9945 18751 9948
rect 18693 9939 18751 9945
rect 19058 9936 19064 9948
rect 19116 9976 19122 9988
rect 19444 9985 19472 10016
rect 19705 10013 19717 10016
rect 19751 10013 19763 10047
rect 19705 10007 19763 10013
rect 19889 10047 19947 10053
rect 19889 10013 19901 10047
rect 19935 10013 19947 10047
rect 19889 10007 19947 10013
rect 19245 9979 19303 9985
rect 19245 9976 19257 9979
rect 19116 9948 19257 9976
rect 19116 9936 19122 9948
rect 19245 9945 19257 9948
rect 19291 9945 19303 9979
rect 19245 9939 19303 9945
rect 19429 9979 19487 9985
rect 19429 9945 19441 9979
rect 19475 9945 19487 9979
rect 19429 9939 19487 9945
rect 19610 9936 19616 9988
rect 19668 9936 19674 9988
rect 19720 9976 19748 10007
rect 20162 10004 20168 10056
rect 20220 10004 20226 10056
rect 20346 10004 20352 10056
rect 20404 10044 20410 10056
rect 20530 10044 20536 10056
rect 20404 10016 20536 10044
rect 20404 10004 20410 10016
rect 20530 10004 20536 10016
rect 20588 10004 20594 10056
rect 24026 10004 24032 10056
rect 24084 10044 24090 10056
rect 24412 10053 24440 10152
rect 24946 10140 24952 10192
rect 25004 10180 25010 10192
rect 25004 10152 25176 10180
rect 25004 10140 25010 10152
rect 24670 10072 24676 10124
rect 24728 10112 24734 10124
rect 25041 10115 25099 10121
rect 25041 10112 25053 10115
rect 24728 10084 25053 10112
rect 24728 10072 24734 10084
rect 25041 10081 25053 10084
rect 25087 10081 25099 10115
rect 25148 10112 25176 10152
rect 25317 10115 25375 10121
rect 25317 10112 25329 10115
rect 25148 10084 25329 10112
rect 25041 10075 25099 10081
rect 25317 10081 25329 10084
rect 25363 10081 25375 10115
rect 25317 10075 25375 10081
rect 24397 10047 24455 10053
rect 24397 10044 24409 10047
rect 24084 10016 24409 10044
rect 24084 10004 24090 10016
rect 24397 10013 24409 10016
rect 24443 10013 24455 10047
rect 24397 10007 24455 10013
rect 24578 10004 24584 10056
rect 24636 10004 24642 10056
rect 20441 9979 20499 9985
rect 19720 9948 20300 9976
rect 19794 9908 19800 9920
rect 16960 9880 19800 9908
rect 19794 9868 19800 9880
rect 19852 9868 19858 9920
rect 20272 9917 20300 9948
rect 20441 9945 20453 9979
rect 20487 9976 20499 9979
rect 20806 9976 20812 9988
rect 20487 9948 20812 9976
rect 20487 9945 20499 9948
rect 20441 9939 20499 9945
rect 20806 9936 20812 9948
rect 20864 9936 20870 9988
rect 21450 9936 21456 9988
rect 21508 9936 21514 9988
rect 23566 9936 23572 9988
rect 23624 9976 23630 9988
rect 24688 9976 24716 10072
rect 24949 10047 25007 10053
rect 24949 10013 24961 10047
rect 24995 10013 25007 10047
rect 24949 10007 25007 10013
rect 23624 9948 24716 9976
rect 23624 9936 23630 9948
rect 20257 9911 20315 9917
rect 20257 9877 20269 9911
rect 20303 9908 20315 9911
rect 20714 9908 20720 9920
rect 20303 9880 20720 9908
rect 20303 9877 20315 9880
rect 20257 9871 20315 9877
rect 20714 9868 20720 9880
rect 20772 9868 20778 9920
rect 20824 9908 20852 9936
rect 22281 9911 22339 9917
rect 22281 9908 22293 9911
rect 20824 9880 22293 9908
rect 22281 9877 22293 9880
rect 22327 9877 22339 9911
rect 24964 9908 24992 10007
rect 25038 9936 25044 9988
rect 25096 9976 25102 9988
rect 25096 9948 25806 9976
rect 25096 9936 25102 9948
rect 25130 9908 25136 9920
rect 24964 9880 25136 9908
rect 22281 9871 22339 9877
rect 25130 9868 25136 9880
rect 25188 9908 25194 9920
rect 26789 9911 26847 9917
rect 26789 9908 26801 9911
rect 25188 9880 26801 9908
rect 25188 9868 25194 9880
rect 26789 9877 26801 9880
rect 26835 9877 26847 9911
rect 26789 9871 26847 9877
rect 1104 9818 28152 9840
rect 1104 9766 4874 9818
rect 4926 9766 4938 9818
rect 4990 9766 5002 9818
rect 5054 9766 5066 9818
rect 5118 9766 5130 9818
rect 5182 9766 28152 9818
rect 1104 9744 28152 9766
rect 9125 9707 9183 9713
rect 9125 9673 9137 9707
rect 9171 9704 9183 9707
rect 9582 9704 9588 9716
rect 9171 9676 9588 9704
rect 9171 9673 9183 9676
rect 9125 9667 9183 9673
rect 9582 9664 9588 9676
rect 9640 9664 9646 9716
rect 11146 9664 11152 9716
rect 11204 9704 11210 9716
rect 18509 9707 18567 9713
rect 11204 9676 17908 9704
rect 11204 9664 11210 9676
rect 8757 9639 8815 9645
rect 8757 9605 8769 9639
rect 8803 9636 8815 9639
rect 8846 9636 8852 9648
rect 8803 9608 8852 9636
rect 8803 9605 8815 9608
rect 8757 9599 8815 9605
rect 8846 9596 8852 9608
rect 8904 9596 8910 9648
rect 8973 9639 9031 9645
rect 8973 9605 8985 9639
rect 9019 9636 9031 9639
rect 9490 9636 9496 9648
rect 9019 9608 9496 9636
rect 9019 9605 9031 9608
rect 8973 9599 9031 9605
rect 9490 9596 9496 9608
rect 9548 9596 9554 9648
rect 13722 9636 13728 9648
rect 13372 9608 13728 9636
rect 12158 9528 12164 9580
rect 12216 9528 12222 9580
rect 12250 9528 12256 9580
rect 12308 9528 12314 9580
rect 12396 9571 12454 9577
rect 12396 9537 12408 9571
rect 12442 9537 12454 9571
rect 12396 9531 12454 9537
rect 12529 9574 12587 9577
rect 12618 9574 12624 9580
rect 12529 9571 12624 9574
rect 12529 9537 12541 9571
rect 12575 9546 12624 9571
rect 12575 9537 12587 9546
rect 12529 9531 12587 9537
rect 12406 9432 12434 9531
rect 12618 9528 12624 9546
rect 12676 9528 12682 9580
rect 12897 9571 12955 9577
rect 12897 9537 12909 9571
rect 12943 9537 12955 9571
rect 12897 9531 12955 9537
rect 12912 9500 12940 9531
rect 12986 9528 12992 9580
rect 13044 9568 13050 9580
rect 13372 9577 13400 9608
rect 13722 9596 13728 9608
rect 13780 9596 13786 9648
rect 13081 9571 13139 9577
rect 13081 9568 13093 9571
rect 13044 9540 13093 9568
rect 13044 9528 13050 9540
rect 13081 9537 13093 9540
rect 13127 9537 13139 9571
rect 13081 9531 13139 9537
rect 13357 9571 13415 9577
rect 13357 9537 13369 9571
rect 13403 9537 13415 9571
rect 13357 9531 13415 9537
rect 13446 9528 13452 9580
rect 13504 9528 13510 9580
rect 13538 9528 13544 9580
rect 13596 9568 13602 9580
rect 13633 9571 13691 9577
rect 13633 9568 13645 9571
rect 13596 9540 13645 9568
rect 13596 9528 13602 9540
rect 13633 9537 13645 9540
rect 13679 9537 13691 9571
rect 13633 9531 13691 9537
rect 12912 9472 13676 9500
rect 12912 9444 12940 9472
rect 13648 9444 13676 9472
rect 12710 9432 12716 9444
rect 12406 9404 12716 9432
rect 12710 9392 12716 9404
rect 12768 9392 12774 9444
rect 12894 9392 12900 9444
rect 12952 9392 12958 9444
rect 12989 9435 13047 9441
rect 12989 9401 13001 9435
rect 13035 9432 13047 9435
rect 13449 9435 13507 9441
rect 13449 9432 13461 9435
rect 13035 9404 13461 9432
rect 13035 9401 13047 9404
rect 12989 9395 13047 9401
rect 13449 9401 13461 9404
rect 13495 9401 13507 9435
rect 13449 9395 13507 9401
rect 13630 9392 13636 9444
rect 13688 9392 13694 9444
rect 17880 9376 17908 9676
rect 18509 9673 18521 9707
rect 18555 9704 18567 9707
rect 18782 9704 18788 9716
rect 18555 9676 18788 9704
rect 18555 9673 18567 9676
rect 18509 9667 18567 9673
rect 18782 9664 18788 9676
rect 18840 9664 18846 9716
rect 21450 9664 21456 9716
rect 21508 9704 21514 9716
rect 21508 9676 21772 9704
rect 21508 9664 21514 9676
rect 18877 9639 18935 9645
rect 18877 9605 18889 9639
rect 18923 9636 18935 9639
rect 19058 9636 19064 9648
rect 18923 9608 19064 9636
rect 18923 9605 18935 9608
rect 18877 9599 18935 9605
rect 19058 9596 19064 9608
rect 19116 9596 19122 9648
rect 20806 9596 20812 9648
rect 20864 9636 20870 9648
rect 20901 9639 20959 9645
rect 20901 9636 20913 9639
rect 20864 9608 20913 9636
rect 20864 9596 20870 9608
rect 20901 9605 20913 9608
rect 20947 9605 20959 9639
rect 21101 9639 21159 9645
rect 21101 9636 21113 9639
rect 20901 9599 20959 9605
rect 21008 9608 21113 9636
rect 18138 9528 18144 9580
rect 18196 9528 18202 9580
rect 18693 9571 18751 9577
rect 18693 9537 18705 9571
rect 18739 9537 18751 9571
rect 18969 9571 19027 9577
rect 18969 9568 18981 9571
rect 18693 9531 18751 9537
rect 18892 9540 18981 9568
rect 18230 9460 18236 9512
rect 18288 9500 18294 9512
rect 18708 9500 18736 9531
rect 18892 9512 18920 9540
rect 18969 9537 18981 9540
rect 19015 9537 19027 9571
rect 18969 9531 19027 9537
rect 20162 9528 20168 9580
rect 20220 9568 20226 9580
rect 21008 9568 21036 9608
rect 21101 9605 21113 9608
rect 21147 9605 21159 9639
rect 21744 9636 21772 9676
rect 21818 9664 21824 9716
rect 21876 9664 21882 9716
rect 25038 9704 25044 9716
rect 21928 9676 25044 9704
rect 21928 9636 21956 9676
rect 25038 9664 25044 9676
rect 25096 9664 25102 9716
rect 22278 9636 22284 9648
rect 21744 9608 21956 9636
rect 22112 9608 22284 9636
rect 21101 9599 21159 9605
rect 22112 9577 22140 9608
rect 22278 9596 22284 9608
rect 22336 9596 22342 9648
rect 20220 9540 21036 9568
rect 22097 9571 22155 9577
rect 20220 9528 20226 9540
rect 22097 9537 22109 9571
rect 22143 9537 22155 9571
rect 22097 9531 22155 9537
rect 22186 9528 22192 9580
rect 22244 9528 22250 9580
rect 22554 9528 22560 9580
rect 22612 9528 22618 9580
rect 24026 9528 24032 9580
rect 24084 9528 24090 9580
rect 24213 9571 24271 9577
rect 24213 9537 24225 9571
rect 24259 9568 24271 9571
rect 24578 9568 24584 9580
rect 24259 9540 24584 9568
rect 24259 9537 24271 9540
rect 24213 9531 24271 9537
rect 24578 9528 24584 9540
rect 24636 9528 24642 9580
rect 18288 9472 18736 9500
rect 18288 9460 18294 9472
rect 18874 9460 18880 9512
rect 18932 9460 18938 9512
rect 22370 9460 22376 9512
rect 22428 9460 22434 9512
rect 18966 9392 18972 9444
rect 19024 9392 19030 9444
rect 21269 9435 21327 9441
rect 21269 9401 21281 9435
rect 21315 9432 21327 9435
rect 22002 9432 22008 9444
rect 21315 9404 22008 9432
rect 21315 9401 21327 9404
rect 21269 9395 21327 9401
rect 22002 9392 22008 9404
rect 22060 9432 22066 9444
rect 22281 9435 22339 9441
rect 22281 9432 22293 9435
rect 22060 9404 22293 9432
rect 22060 9392 22066 9404
rect 22281 9401 22293 9404
rect 22327 9401 22339 9435
rect 22281 9395 22339 9401
rect 8938 9324 8944 9376
rect 8996 9324 9002 9376
rect 11977 9367 12035 9373
rect 11977 9333 11989 9367
rect 12023 9364 12035 9367
rect 12250 9364 12256 9376
rect 12023 9336 12256 9364
rect 12023 9333 12035 9336
rect 11977 9327 12035 9333
rect 12250 9324 12256 9336
rect 12308 9324 12314 9376
rect 12342 9324 12348 9376
rect 12400 9364 12406 9376
rect 12621 9367 12679 9373
rect 12621 9364 12633 9367
rect 12400 9336 12633 9364
rect 12400 9324 12406 9336
rect 12621 9333 12633 9336
rect 12667 9333 12679 9367
rect 12621 9327 12679 9333
rect 13173 9367 13231 9373
rect 13173 9333 13185 9367
rect 13219 9364 13231 9367
rect 13262 9364 13268 9376
rect 13219 9336 13268 9364
rect 13219 9333 13231 9336
rect 13173 9327 13231 9333
rect 13262 9324 13268 9336
rect 13320 9324 13326 9376
rect 17862 9324 17868 9376
rect 17920 9364 17926 9376
rect 19610 9364 19616 9376
rect 17920 9336 19616 9364
rect 17920 9324 17926 9336
rect 19610 9324 19616 9336
rect 19668 9364 19674 9376
rect 19978 9364 19984 9376
rect 19668 9336 19984 9364
rect 19668 9324 19674 9336
rect 19978 9324 19984 9336
rect 20036 9324 20042 9376
rect 20714 9324 20720 9376
rect 20772 9364 20778 9376
rect 21082 9364 21088 9376
rect 20772 9336 21088 9364
rect 20772 9324 20778 9336
rect 21082 9324 21088 9336
rect 21140 9324 21146 9376
rect 23658 9324 23664 9376
rect 23716 9364 23722 9376
rect 24213 9367 24271 9373
rect 24213 9364 24225 9367
rect 23716 9336 24225 9364
rect 23716 9324 23722 9336
rect 24213 9333 24225 9336
rect 24259 9333 24271 9367
rect 24213 9327 24271 9333
rect 24489 9367 24547 9373
rect 24489 9333 24501 9367
rect 24535 9364 24547 9367
rect 24854 9364 24860 9376
rect 24535 9336 24860 9364
rect 24535 9333 24547 9336
rect 24489 9327 24547 9333
rect 24854 9324 24860 9336
rect 24912 9324 24918 9376
rect 1104 9274 28152 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 28152 9274
rect 1104 9200 28152 9222
rect 6270 9120 6276 9172
rect 6328 9120 6334 9172
rect 8205 9163 8263 9169
rect 8205 9129 8217 9163
rect 8251 9160 8263 9163
rect 8938 9160 8944 9172
rect 8251 9132 8944 9160
rect 8251 9129 8263 9132
rect 8205 9123 8263 9129
rect 8938 9120 8944 9132
rect 8996 9120 9002 9172
rect 11698 9120 11704 9172
rect 11756 9160 11762 9172
rect 11885 9163 11943 9169
rect 11885 9160 11897 9163
rect 11756 9132 11897 9160
rect 11756 9120 11762 9132
rect 11885 9129 11897 9132
rect 11931 9160 11943 9163
rect 11931 9132 12434 9160
rect 11931 9129 11943 9132
rect 11885 9123 11943 9129
rect 4798 8984 4804 9036
rect 4856 9024 4862 9036
rect 4985 9027 5043 9033
rect 4985 9024 4997 9027
rect 4856 8996 4997 9024
rect 4856 8984 4862 8996
rect 4985 8993 4997 8996
rect 5031 8993 5043 9027
rect 4985 8987 5043 8993
rect 5626 8984 5632 9036
rect 5684 9024 5690 9036
rect 9953 9027 10011 9033
rect 5684 8996 6132 9024
rect 5684 8984 5690 8996
rect 6104 8968 6132 8996
rect 9953 8993 9965 9027
rect 9999 9024 10011 9027
rect 10594 9024 10600 9036
rect 9999 8996 10600 9024
rect 9999 8993 10011 8996
rect 9953 8987 10011 8993
rect 10594 8984 10600 8996
rect 10652 8984 10658 9036
rect 12406 9024 12434 9132
rect 12802 9120 12808 9172
rect 12860 9160 12866 9172
rect 13081 9163 13139 9169
rect 13081 9160 13093 9163
rect 12860 9132 13093 9160
rect 12860 9120 12866 9132
rect 13081 9129 13093 9132
rect 13127 9129 13139 9163
rect 13081 9123 13139 9129
rect 16574 9120 16580 9172
rect 16632 9160 16638 9172
rect 16853 9163 16911 9169
rect 16853 9160 16865 9163
rect 16632 9132 16865 9160
rect 16632 9120 16638 9132
rect 16853 9129 16865 9132
rect 16899 9129 16911 9163
rect 18230 9160 18236 9172
rect 16853 9123 16911 9129
rect 17236 9132 18236 9160
rect 12618 9052 12624 9104
rect 12676 9092 12682 9104
rect 12986 9092 12992 9104
rect 12676 9064 12992 9092
rect 12676 9052 12682 9064
rect 12986 9052 12992 9064
rect 13044 9052 13050 9104
rect 17236 9092 17264 9132
rect 18230 9120 18236 9132
rect 18288 9120 18294 9172
rect 23382 9120 23388 9172
rect 23440 9120 23446 9172
rect 24857 9163 24915 9169
rect 24857 9129 24869 9163
rect 24903 9160 24915 9163
rect 25130 9160 25136 9172
rect 24903 9132 25136 9160
rect 24903 9129 24915 9132
rect 24857 9123 24915 9129
rect 25130 9120 25136 9132
rect 25188 9120 25194 9172
rect 16132 9064 17264 9092
rect 12406 8996 12480 9024
rect 5077 8959 5135 8965
rect 5077 8925 5089 8959
rect 5123 8956 5135 8959
rect 5350 8956 5356 8968
rect 5123 8928 5356 8956
rect 5123 8925 5135 8928
rect 5077 8919 5135 8925
rect 5350 8916 5356 8928
rect 5408 8916 5414 8968
rect 5810 8916 5816 8968
rect 5868 8916 5874 8968
rect 5902 8916 5908 8968
rect 5960 8916 5966 8968
rect 5997 8959 6055 8965
rect 5997 8925 6009 8959
rect 6043 8925 6055 8959
rect 5997 8919 6055 8925
rect 6012 8888 6040 8919
rect 6086 8916 6092 8968
rect 6144 8916 6150 8968
rect 8110 8916 8116 8968
rect 8168 8916 8174 8968
rect 8297 8959 8355 8965
rect 8297 8925 8309 8959
rect 8343 8925 8355 8959
rect 8297 8919 8355 8925
rect 6178 8888 6184 8900
rect 6012 8860 6184 8888
rect 6178 8848 6184 8860
rect 6236 8848 6242 8900
rect 8018 8848 8024 8900
rect 8076 8888 8082 8900
rect 8312 8888 8340 8919
rect 9674 8916 9680 8968
rect 9732 8916 9738 8968
rect 9769 8959 9827 8965
rect 9769 8925 9781 8959
rect 9815 8925 9827 8959
rect 9769 8919 9827 8925
rect 8076 8860 8340 8888
rect 8076 8848 8082 8860
rect 9582 8848 9588 8900
rect 9640 8888 9646 8900
rect 9784 8888 9812 8919
rect 9640 8860 9812 8888
rect 10612 8888 10640 8984
rect 12066 8916 12072 8968
rect 12124 8916 12130 8968
rect 12250 8916 12256 8968
rect 12308 8916 12314 8968
rect 12342 8916 12348 8968
rect 12400 8916 12406 8968
rect 12452 8965 12480 8996
rect 12437 8959 12495 8965
rect 12437 8925 12449 8959
rect 12483 8925 12495 8959
rect 12437 8919 12495 8925
rect 13078 8916 13084 8968
rect 13136 8916 13142 8968
rect 13265 8959 13323 8965
rect 13265 8925 13277 8959
rect 13311 8956 13323 8959
rect 14090 8956 14096 8968
rect 13311 8928 14096 8956
rect 13311 8925 13323 8928
rect 13265 8919 13323 8925
rect 14090 8916 14096 8928
rect 14148 8916 14154 8968
rect 16132 8888 16160 9064
rect 17310 9052 17316 9104
rect 17368 9092 17374 9104
rect 17405 9095 17463 9101
rect 17405 9092 17417 9095
rect 17368 9064 17417 9092
rect 17368 9052 17374 9064
rect 17405 9061 17417 9064
rect 17451 9061 17463 9095
rect 24949 9095 25007 9101
rect 24949 9092 24961 9095
rect 17405 9055 17463 9061
rect 23492 9064 24961 9092
rect 16574 8984 16580 9036
rect 16632 9024 16638 9036
rect 16632 8996 17264 9024
rect 16632 8984 16638 8996
rect 16206 8916 16212 8968
rect 16264 8956 16270 8968
rect 17236 8965 17264 8996
rect 23382 8984 23388 9036
rect 23440 9024 23446 9036
rect 23492 9024 23520 9064
rect 24949 9061 24961 9064
rect 24995 9061 25007 9095
rect 24949 9055 25007 9061
rect 24121 9027 24179 9033
rect 24121 9024 24133 9027
rect 23440 8996 23520 9024
rect 23584 8996 24133 9024
rect 23440 8984 23446 8996
rect 23584 8965 23612 8996
rect 24121 8993 24133 8996
rect 24167 8993 24179 9027
rect 24121 8987 24179 8993
rect 24762 8984 24768 9036
rect 24820 8984 24826 9036
rect 17129 8959 17187 8965
rect 17129 8956 17141 8959
rect 16264 8928 17141 8956
rect 16264 8916 16270 8928
rect 16868 8897 16896 8928
rect 17129 8925 17141 8928
rect 17175 8925 17187 8959
rect 17129 8919 17187 8925
rect 17221 8959 17279 8965
rect 17221 8925 17233 8959
rect 17267 8925 17279 8959
rect 17221 8919 17279 8925
rect 23017 8959 23075 8965
rect 23017 8925 23029 8959
rect 23063 8925 23075 8959
rect 23017 8919 23075 8925
rect 23109 8959 23167 8965
rect 23109 8925 23121 8959
rect 23155 8956 23167 8959
rect 23569 8959 23627 8965
rect 23569 8956 23581 8959
rect 23155 8928 23581 8956
rect 23155 8925 23167 8928
rect 23109 8919 23167 8925
rect 23569 8925 23581 8928
rect 23615 8925 23627 8959
rect 23569 8919 23627 8925
rect 10612 8860 16160 8888
rect 16669 8891 16727 8897
rect 9640 8848 9646 8860
rect 16669 8857 16681 8891
rect 16715 8857 16727 8891
rect 16868 8891 16927 8897
rect 16868 8860 16881 8891
rect 16669 8851 16727 8857
rect 16869 8857 16881 8860
rect 16915 8857 16927 8891
rect 17405 8891 17463 8897
rect 17405 8888 17417 8891
rect 16869 8851 16927 8857
rect 16960 8860 17417 8888
rect 5445 8823 5503 8829
rect 5445 8789 5457 8823
rect 5491 8820 5503 8823
rect 5902 8820 5908 8832
rect 5491 8792 5908 8820
rect 5491 8789 5503 8792
rect 5445 8783 5503 8789
rect 5902 8780 5908 8792
rect 5960 8780 5966 8832
rect 6196 8820 6224 8848
rect 11698 8820 11704 8832
rect 6196 8792 11704 8820
rect 11698 8780 11704 8792
rect 11756 8780 11762 8832
rect 12434 8780 12440 8832
rect 12492 8820 12498 8832
rect 12529 8823 12587 8829
rect 12529 8820 12541 8823
rect 12492 8792 12541 8820
rect 12492 8780 12498 8792
rect 12529 8789 12541 8792
rect 12575 8789 12587 8823
rect 16684 8820 16712 8851
rect 16960 8820 16988 8860
rect 17405 8857 17417 8860
rect 17451 8888 17463 8891
rect 17954 8888 17960 8900
rect 17451 8860 17960 8888
rect 17451 8857 17463 8860
rect 17405 8851 17463 8857
rect 17954 8848 17960 8860
rect 18012 8848 18018 8900
rect 23032 8888 23060 8919
rect 23658 8916 23664 8968
rect 23716 8916 23722 8968
rect 23937 8959 23995 8965
rect 23937 8925 23949 8959
rect 23983 8925 23995 8959
rect 23937 8919 23995 8925
rect 23676 8888 23704 8916
rect 23032 8860 23704 8888
rect 23750 8848 23756 8900
rect 23808 8848 23814 8900
rect 23952 8888 23980 8919
rect 24026 8916 24032 8968
rect 24084 8916 24090 8968
rect 24210 8916 24216 8968
rect 24268 8916 24274 8968
rect 24581 8959 24639 8965
rect 24581 8925 24593 8959
rect 24627 8925 24639 8959
rect 24581 8919 24639 8925
rect 24118 8888 24124 8900
rect 23952 8860 24124 8888
rect 24118 8848 24124 8860
rect 24176 8848 24182 8900
rect 16684 8792 16988 8820
rect 17037 8823 17095 8829
rect 12529 8783 12587 8789
rect 17037 8789 17049 8823
rect 17083 8820 17095 8823
rect 17126 8820 17132 8832
rect 17083 8792 17132 8820
rect 17083 8789 17095 8792
rect 17037 8783 17095 8789
rect 17126 8780 17132 8792
rect 17184 8780 17190 8832
rect 17586 8780 17592 8832
rect 17644 8820 17650 8832
rect 18414 8820 18420 8832
rect 17644 8792 18420 8820
rect 17644 8780 17650 8792
rect 18414 8780 18420 8792
rect 18472 8820 18478 8832
rect 18782 8820 18788 8832
rect 18472 8792 18788 8820
rect 18472 8780 18478 8792
rect 18782 8780 18788 8792
rect 18840 8780 18846 8832
rect 23293 8823 23351 8829
rect 23293 8789 23305 8823
rect 23339 8820 23351 8823
rect 23934 8820 23940 8832
rect 23339 8792 23940 8820
rect 23339 8789 23351 8792
rect 23293 8783 23351 8789
rect 23934 8780 23940 8792
rect 23992 8780 23998 8832
rect 24210 8780 24216 8832
rect 24268 8820 24274 8832
rect 24397 8823 24455 8829
rect 24397 8820 24409 8823
rect 24268 8792 24409 8820
rect 24268 8780 24274 8792
rect 24397 8789 24409 8792
rect 24443 8789 24455 8823
rect 24596 8820 24624 8919
rect 24854 8916 24860 8968
rect 24912 8916 24918 8968
rect 24872 8888 24900 8916
rect 25101 8891 25159 8897
rect 25101 8888 25113 8891
rect 24872 8860 25113 8888
rect 25101 8857 25113 8860
rect 25147 8857 25159 8891
rect 25101 8851 25159 8857
rect 25317 8891 25375 8897
rect 25317 8857 25329 8891
rect 25363 8857 25375 8891
rect 25317 8851 25375 8857
rect 24946 8820 24952 8832
rect 24596 8792 24952 8820
rect 24397 8783 24455 8789
rect 24946 8780 24952 8792
rect 25004 8820 25010 8832
rect 25332 8820 25360 8851
rect 25004 8792 25360 8820
rect 25004 8780 25010 8792
rect 1104 8730 28152 8752
rect 1104 8678 4874 8730
rect 4926 8678 4938 8730
rect 4990 8678 5002 8730
rect 5054 8678 5066 8730
rect 5118 8678 5130 8730
rect 5182 8678 28152 8730
rect 1104 8656 28152 8678
rect 5353 8619 5411 8625
rect 5353 8585 5365 8619
rect 5399 8616 5411 8619
rect 5810 8616 5816 8628
rect 5399 8588 5816 8616
rect 5399 8585 5411 8588
rect 5353 8579 5411 8585
rect 5810 8576 5816 8588
rect 5868 8576 5874 8628
rect 9674 8576 9680 8628
rect 9732 8576 9738 8628
rect 11698 8576 11704 8628
rect 11756 8576 11762 8628
rect 14185 8619 14243 8625
rect 14185 8585 14197 8619
rect 14231 8616 14243 8619
rect 14366 8616 14372 8628
rect 14231 8588 14372 8616
rect 14231 8585 14243 8588
rect 14185 8579 14243 8585
rect 14366 8576 14372 8588
rect 14424 8576 14430 8628
rect 24210 8616 24216 8628
rect 14752 8588 24216 8616
rect 6089 8551 6147 8557
rect 6089 8517 6101 8551
rect 6135 8548 6147 8551
rect 9493 8551 9551 8557
rect 9493 8548 9505 8551
rect 6135 8520 6592 8548
rect 6135 8517 6147 8520
rect 6089 8511 6147 8517
rect 4798 8440 4804 8492
rect 4856 8480 4862 8492
rect 5169 8483 5227 8489
rect 5169 8480 5181 8483
rect 4856 8452 5181 8480
rect 4856 8440 4862 8452
rect 5169 8449 5181 8452
rect 5215 8449 5227 8483
rect 5169 8443 5227 8449
rect 5350 8440 5356 8492
rect 5408 8440 5414 8492
rect 5534 8440 5540 8492
rect 5592 8440 5598 8492
rect 5810 8440 5816 8492
rect 5868 8480 5874 8492
rect 5994 8480 6000 8492
rect 5868 8452 6000 8480
rect 5868 8440 5874 8452
rect 5994 8440 6000 8452
rect 6052 8440 6058 8492
rect 6178 8440 6184 8492
rect 6236 8440 6242 8492
rect 6564 8489 6592 8520
rect 8404 8520 9505 8548
rect 6549 8483 6607 8489
rect 6549 8449 6561 8483
rect 6595 8449 6607 8483
rect 6549 8443 6607 8449
rect 8018 8440 8024 8492
rect 8076 8440 8082 8492
rect 5902 8372 5908 8424
rect 5960 8412 5966 8424
rect 6457 8415 6515 8421
rect 6457 8412 6469 8415
rect 5960 8384 6469 8412
rect 5960 8372 5966 8384
rect 6457 8381 6469 8384
rect 6503 8381 6515 8415
rect 6457 8375 6515 8381
rect 7929 8415 7987 8421
rect 7929 8381 7941 8415
rect 7975 8412 7987 8415
rect 8110 8412 8116 8424
rect 7975 8384 8116 8412
rect 7975 8381 7987 8384
rect 7929 8375 7987 8381
rect 6917 8347 6975 8353
rect 6917 8313 6929 8347
rect 6963 8344 6975 8347
rect 7944 8344 7972 8375
rect 8110 8372 8116 8384
rect 8168 8372 8174 8424
rect 8404 8421 8432 8520
rect 9493 8517 9505 8520
rect 9539 8517 9551 8551
rect 9493 8511 9551 8517
rect 9309 8483 9367 8489
rect 9309 8449 9321 8483
rect 9355 8449 9367 8483
rect 9508 8480 9536 8511
rect 9582 8508 9588 8560
rect 9640 8548 9646 8560
rect 9861 8551 9919 8557
rect 9861 8548 9873 8551
rect 9640 8520 9873 8548
rect 9640 8508 9646 8520
rect 9861 8517 9873 8520
rect 9907 8517 9919 8551
rect 9861 8511 9919 8517
rect 12713 8551 12771 8557
rect 12713 8517 12725 8551
rect 12759 8548 12771 8551
rect 13078 8548 13084 8560
rect 12759 8520 13084 8548
rect 12759 8517 12771 8520
rect 12713 8511 12771 8517
rect 13078 8508 13084 8520
rect 13136 8548 13142 8560
rect 13136 8520 14688 8548
rect 13136 8508 13142 8520
rect 9769 8483 9827 8489
rect 9769 8480 9781 8483
rect 9508 8452 9781 8480
rect 9309 8443 9367 8449
rect 9769 8449 9781 8452
rect 9815 8449 9827 8483
rect 9769 8443 9827 8449
rect 8389 8415 8447 8421
rect 8389 8381 8401 8415
rect 8435 8381 8447 8415
rect 8389 8375 8447 8381
rect 6963 8316 7972 8344
rect 9324 8344 9352 8443
rect 9950 8440 9956 8492
rect 10008 8440 10014 8492
rect 11609 8483 11667 8489
rect 11609 8449 11621 8483
rect 11655 8480 11667 8483
rect 12621 8483 12679 8489
rect 12621 8480 12633 8483
rect 11655 8452 12633 8480
rect 11655 8449 11667 8452
rect 11609 8443 11667 8449
rect 12621 8449 12633 8452
rect 12667 8449 12679 8483
rect 12621 8443 12679 8449
rect 9582 8372 9588 8424
rect 9640 8412 9646 8424
rect 11624 8412 11652 8443
rect 12802 8440 12808 8492
rect 12860 8440 12866 8492
rect 13906 8440 13912 8492
rect 13964 8480 13970 8492
rect 14660 8489 14688 8520
rect 14752 8489 14780 8588
rect 24210 8576 24216 8588
rect 24268 8576 24274 8628
rect 24854 8576 24860 8628
rect 24912 8616 24918 8628
rect 25409 8619 25467 8625
rect 25409 8616 25421 8619
rect 24912 8588 25421 8616
rect 24912 8576 24918 8588
rect 25409 8585 25421 8588
rect 25455 8585 25467 8619
rect 25409 8579 25467 8585
rect 17310 8508 17316 8560
rect 17368 8508 17374 8560
rect 18892 8520 19656 8548
rect 14369 8483 14427 8489
rect 14369 8480 14381 8483
rect 13964 8452 14381 8480
rect 13964 8440 13970 8452
rect 14369 8449 14381 8452
rect 14415 8449 14427 8483
rect 14369 8443 14427 8449
rect 14461 8483 14519 8489
rect 14461 8449 14473 8483
rect 14507 8449 14519 8483
rect 14461 8443 14519 8449
rect 14645 8483 14703 8489
rect 14645 8449 14657 8483
rect 14691 8449 14703 8483
rect 14645 8443 14703 8449
rect 14737 8483 14795 8489
rect 14737 8449 14749 8483
rect 14783 8449 14795 8483
rect 14737 8443 14795 8449
rect 9640 8384 11652 8412
rect 9640 8372 9646 8384
rect 13814 8372 13820 8424
rect 13872 8412 13878 8424
rect 14476 8412 14504 8443
rect 14918 8440 14924 8492
rect 14976 8480 14982 8492
rect 16850 8480 16856 8492
rect 14976 8452 16856 8480
rect 14976 8440 14982 8452
rect 16850 8440 16856 8452
rect 16908 8480 16914 8492
rect 17037 8483 17095 8489
rect 17037 8480 17049 8483
rect 16908 8452 17049 8480
rect 16908 8440 16914 8452
rect 17037 8449 17049 8452
rect 17083 8449 17095 8483
rect 17037 8443 17095 8449
rect 13872 8384 14504 8412
rect 13872 8372 13878 8384
rect 9950 8344 9956 8356
rect 9324 8316 9956 8344
rect 6963 8313 6975 8316
rect 6917 8307 6975 8313
rect 9950 8304 9956 8316
rect 10008 8304 10014 8356
rect 11624 8316 11836 8344
rect 5629 8279 5687 8285
rect 5629 8245 5641 8279
rect 5675 8276 5687 8279
rect 5810 8276 5816 8288
rect 5675 8248 5816 8276
rect 5675 8245 5687 8248
rect 5629 8239 5687 8245
rect 5810 8236 5816 8248
rect 5868 8236 5874 8288
rect 10870 8236 10876 8288
rect 10928 8276 10934 8288
rect 11624 8276 11652 8316
rect 10928 8248 11652 8276
rect 11808 8276 11836 8316
rect 13446 8304 13452 8356
rect 13504 8344 13510 8356
rect 13722 8344 13728 8356
rect 13504 8316 13728 8344
rect 13504 8304 13510 8316
rect 13722 8304 13728 8316
rect 13780 8344 13786 8356
rect 14918 8344 14924 8356
rect 13780 8316 14924 8344
rect 13780 8304 13786 8316
rect 14918 8304 14924 8316
rect 14976 8304 14982 8356
rect 17052 8344 17080 8443
rect 17126 8440 17132 8492
rect 17184 8480 17190 8492
rect 18892 8480 18920 8520
rect 17184 8452 18920 8480
rect 17184 8440 17190 8452
rect 18966 8440 18972 8492
rect 19024 8480 19030 8492
rect 19628 8489 19656 8520
rect 19978 8508 19984 8560
rect 20036 8548 20042 8560
rect 23201 8551 23259 8557
rect 23201 8548 23213 8551
rect 20036 8520 20208 8548
rect 20036 8508 20042 8520
rect 20180 8489 20208 8520
rect 22066 8520 23213 8548
rect 19429 8483 19487 8489
rect 19429 8480 19441 8483
rect 19024 8452 19441 8480
rect 19024 8440 19030 8452
rect 19429 8449 19441 8452
rect 19475 8449 19487 8483
rect 19429 8443 19487 8449
rect 19613 8483 19671 8489
rect 19613 8449 19625 8483
rect 19659 8480 19671 8483
rect 19889 8483 19947 8489
rect 19889 8480 19901 8483
rect 19659 8452 19901 8480
rect 19659 8449 19671 8452
rect 19613 8443 19671 8449
rect 19889 8449 19901 8452
rect 19935 8449 19947 8483
rect 19889 8443 19947 8449
rect 20073 8483 20131 8489
rect 20073 8449 20085 8483
rect 20119 8449 20131 8483
rect 20073 8443 20131 8449
rect 20165 8483 20223 8489
rect 20165 8449 20177 8483
rect 20211 8449 20223 8483
rect 20165 8443 20223 8449
rect 18138 8372 18144 8424
rect 18196 8412 18202 8424
rect 18506 8412 18512 8424
rect 18196 8384 18512 8412
rect 18196 8372 18202 8384
rect 18506 8372 18512 8384
rect 18564 8412 18570 8424
rect 19061 8415 19119 8421
rect 19061 8412 19073 8415
rect 18564 8384 19073 8412
rect 18564 8372 18570 8384
rect 19061 8381 19073 8384
rect 19107 8381 19119 8415
rect 19444 8412 19472 8443
rect 20088 8412 20116 8443
rect 20898 8440 20904 8492
rect 20956 8480 20962 8492
rect 22066 8480 22094 8520
rect 23201 8517 23213 8520
rect 23247 8517 23259 8551
rect 23201 8511 23259 8517
rect 23382 8508 23388 8560
rect 23440 8508 23446 8560
rect 23934 8508 23940 8560
rect 23992 8508 23998 8560
rect 20956 8452 22094 8480
rect 22741 8483 22799 8489
rect 20956 8440 20962 8452
rect 22741 8449 22753 8483
rect 22787 8480 22799 8483
rect 22787 8452 23244 8480
rect 22787 8449 22799 8452
rect 22741 8443 22799 8449
rect 19444 8384 20116 8412
rect 19061 8375 19119 8381
rect 20254 8372 20260 8424
rect 20312 8412 20318 8424
rect 22002 8412 22008 8424
rect 20312 8384 22008 8412
rect 20312 8372 20318 8384
rect 22002 8372 22008 8384
rect 22060 8372 22066 8424
rect 23216 8412 23244 8452
rect 23290 8440 23296 8492
rect 23348 8440 23354 8492
rect 23566 8440 23572 8492
rect 23624 8480 23630 8492
rect 23661 8483 23719 8489
rect 23661 8480 23673 8483
rect 23624 8452 23673 8480
rect 23624 8440 23630 8452
rect 23661 8449 23673 8452
rect 23707 8449 23719 8483
rect 23661 8443 23719 8449
rect 25038 8440 25044 8492
rect 25096 8440 25102 8492
rect 24026 8412 24032 8424
rect 23216 8384 23428 8412
rect 19426 8344 19432 8356
rect 16684 8316 16988 8344
rect 17052 8316 19432 8344
rect 15930 8276 15936 8288
rect 11808 8248 15936 8276
rect 10928 8236 10934 8248
rect 15930 8236 15936 8248
rect 15988 8236 15994 8288
rect 16114 8236 16120 8288
rect 16172 8276 16178 8288
rect 16684 8276 16712 8316
rect 16172 8248 16712 8276
rect 16172 8236 16178 8248
rect 16758 8236 16764 8288
rect 16816 8276 16822 8288
rect 16853 8279 16911 8285
rect 16853 8276 16865 8279
rect 16816 8248 16865 8276
rect 16816 8236 16822 8248
rect 16853 8245 16865 8248
rect 16899 8245 16911 8279
rect 16960 8276 16988 8316
rect 19426 8304 19432 8316
rect 19484 8304 19490 8356
rect 19702 8304 19708 8356
rect 19760 8344 19766 8356
rect 19797 8347 19855 8353
rect 19797 8344 19809 8347
rect 19760 8316 19809 8344
rect 19760 8304 19766 8316
rect 19797 8313 19809 8316
rect 19843 8344 19855 8347
rect 20162 8344 20168 8356
rect 19843 8316 20168 8344
rect 19843 8313 19855 8316
rect 19797 8307 19855 8313
rect 20162 8304 20168 8316
rect 20220 8304 20226 8356
rect 22922 8344 22928 8356
rect 22066 8316 22928 8344
rect 17313 8279 17371 8285
rect 17313 8276 17325 8279
rect 16960 8248 17325 8276
rect 16853 8239 16911 8245
rect 17313 8245 17325 8248
rect 17359 8276 17371 8279
rect 19518 8276 19524 8288
rect 17359 8248 19524 8276
rect 17359 8245 17371 8248
rect 17313 8239 17371 8245
rect 19518 8236 19524 8248
rect 19576 8236 19582 8288
rect 19886 8236 19892 8288
rect 19944 8236 19950 8288
rect 20257 8279 20315 8285
rect 20257 8245 20269 8279
rect 20303 8276 20315 8279
rect 20622 8276 20628 8288
rect 20303 8248 20628 8276
rect 20303 8245 20315 8248
rect 20257 8239 20315 8245
rect 20622 8236 20628 8248
rect 20680 8236 20686 8288
rect 20990 8236 20996 8288
rect 21048 8276 21054 8288
rect 21174 8276 21180 8288
rect 21048 8248 21180 8276
rect 21048 8236 21054 8248
rect 21174 8236 21180 8248
rect 21232 8276 21238 8288
rect 22066 8276 22094 8316
rect 22922 8304 22928 8316
rect 22980 8304 22986 8356
rect 23017 8347 23075 8353
rect 23017 8313 23029 8347
rect 23063 8313 23075 8347
rect 23017 8307 23075 8313
rect 21232 8248 22094 8276
rect 21232 8236 21238 8248
rect 22278 8236 22284 8288
rect 22336 8276 22342 8288
rect 22833 8279 22891 8285
rect 22833 8276 22845 8279
rect 22336 8248 22845 8276
rect 22336 8236 22342 8248
rect 22833 8245 22845 8248
rect 22879 8276 22891 8279
rect 23032 8276 23060 8307
rect 22879 8248 23060 8276
rect 23400 8276 23428 8384
rect 23584 8384 24032 8412
rect 23474 8304 23480 8356
rect 23532 8344 23538 8356
rect 23584 8353 23612 8384
rect 24026 8372 24032 8384
rect 24084 8372 24090 8424
rect 23569 8347 23627 8353
rect 23569 8344 23581 8347
rect 23532 8316 23581 8344
rect 23532 8304 23538 8316
rect 23569 8313 23581 8316
rect 23615 8313 23627 8347
rect 23569 8307 23627 8313
rect 24302 8276 24308 8288
rect 23400 8248 24308 8276
rect 22879 8245 22891 8248
rect 22833 8239 22891 8245
rect 24302 8236 24308 8248
rect 24360 8236 24366 8288
rect 1104 8186 28152 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 28152 8186
rect 1104 8112 28152 8134
rect 5261 8075 5319 8081
rect 5261 8041 5273 8075
rect 5307 8072 5319 8075
rect 5350 8072 5356 8084
rect 5307 8044 5356 8072
rect 5307 8041 5319 8044
rect 5261 8035 5319 8041
rect 5350 8032 5356 8044
rect 5408 8032 5414 8084
rect 6181 8075 6239 8081
rect 6181 8041 6193 8075
rect 6227 8072 6239 8075
rect 6546 8072 6552 8084
rect 6227 8044 6552 8072
rect 6227 8041 6239 8044
rect 6181 8035 6239 8041
rect 6196 8004 6224 8035
rect 6546 8032 6552 8044
rect 6604 8072 6610 8084
rect 8478 8072 8484 8084
rect 6604 8044 8484 8072
rect 6604 8032 6610 8044
rect 8478 8032 8484 8044
rect 8536 8072 8542 8084
rect 9582 8072 9588 8084
rect 8536 8044 9588 8072
rect 8536 8032 8542 8044
rect 9582 8032 9588 8044
rect 9640 8032 9646 8084
rect 10781 8075 10839 8081
rect 10781 8041 10793 8075
rect 10827 8072 10839 8075
rect 12618 8072 12624 8084
rect 10827 8044 12624 8072
rect 10827 8041 10839 8044
rect 10781 8035 10839 8041
rect 12618 8032 12624 8044
rect 12676 8032 12682 8084
rect 13170 8032 13176 8084
rect 13228 8032 13234 8084
rect 13541 8075 13599 8081
rect 13541 8041 13553 8075
rect 13587 8072 13599 8075
rect 13906 8072 13912 8084
rect 13587 8044 13912 8072
rect 13587 8041 13599 8044
rect 13541 8035 13599 8041
rect 13906 8032 13912 8044
rect 13964 8032 13970 8084
rect 15933 8075 15991 8081
rect 15933 8041 15945 8075
rect 15979 8072 15991 8075
rect 16761 8075 16819 8081
rect 16761 8072 16773 8075
rect 15979 8044 16773 8072
rect 15979 8041 15991 8044
rect 15933 8035 15991 8041
rect 16761 8041 16773 8044
rect 16807 8041 16819 8075
rect 16761 8035 16819 8041
rect 17218 8032 17224 8084
rect 17276 8032 17282 8084
rect 19613 8075 19671 8081
rect 19613 8041 19625 8075
rect 19659 8072 19671 8075
rect 19886 8072 19892 8084
rect 19659 8044 19892 8072
rect 19659 8041 19671 8044
rect 19613 8035 19671 8041
rect 19886 8032 19892 8044
rect 19944 8032 19950 8084
rect 20070 8032 20076 8084
rect 20128 8032 20134 8084
rect 21177 8075 21235 8081
rect 21177 8041 21189 8075
rect 21223 8041 21235 8075
rect 21177 8035 21235 8041
rect 5552 7976 6224 8004
rect 15841 8007 15899 8013
rect 4614 7936 4620 7948
rect 4356 7908 4620 7936
rect 4356 7877 4384 7908
rect 4614 7896 4620 7908
rect 4672 7936 4678 7948
rect 5552 7945 5580 7976
rect 15841 7973 15853 8007
rect 15887 8004 15899 8007
rect 16022 8004 16028 8016
rect 15887 7976 16028 8004
rect 15887 7973 15899 7976
rect 15841 7967 15899 7973
rect 16022 7964 16028 7976
rect 16080 7964 16086 8016
rect 16942 7964 16948 8016
rect 17000 8004 17006 8016
rect 17000 7976 19380 8004
rect 17000 7964 17006 7976
rect 4709 7939 4767 7945
rect 4709 7936 4721 7939
rect 4672 7908 4721 7936
rect 4672 7896 4678 7908
rect 4709 7905 4721 7908
rect 4755 7905 4767 7939
rect 4709 7899 4767 7905
rect 5169 7939 5227 7945
rect 5169 7905 5181 7939
rect 5215 7905 5227 7939
rect 5169 7899 5227 7905
rect 5537 7939 5595 7945
rect 5537 7905 5549 7939
rect 5583 7905 5595 7939
rect 5537 7899 5595 7905
rect 5629 7939 5687 7945
rect 5629 7905 5641 7939
rect 5675 7936 5687 7939
rect 5810 7936 5816 7948
rect 5675 7908 5816 7936
rect 5675 7905 5687 7908
rect 5629 7899 5687 7905
rect 4341 7871 4399 7877
rect 4341 7837 4353 7871
rect 4387 7837 4399 7871
rect 4341 7831 4399 7837
rect 4525 7871 4583 7877
rect 4525 7837 4537 7871
rect 4571 7868 4583 7871
rect 4798 7868 4804 7880
rect 4571 7840 4804 7868
rect 4571 7837 4583 7840
rect 4525 7831 4583 7837
rect 4798 7828 4804 7840
rect 4856 7828 4862 7880
rect 5184 7868 5212 7899
rect 5810 7896 5816 7908
rect 5868 7896 5874 7948
rect 16853 7939 16911 7945
rect 6288 7908 12664 7936
rect 5442 7868 5448 7880
rect 5184 7840 5448 7868
rect 5442 7828 5448 7840
rect 5500 7828 5506 7880
rect 5721 7871 5779 7877
rect 5721 7837 5733 7871
rect 5767 7837 5779 7871
rect 5721 7831 5779 7837
rect 4433 7803 4491 7809
rect 4433 7769 4445 7803
rect 4479 7800 4491 7803
rect 5736 7800 5764 7831
rect 6086 7828 6092 7880
rect 6144 7868 6150 7880
rect 6288 7877 6316 7908
rect 6273 7871 6331 7877
rect 6273 7868 6285 7871
rect 6144 7840 6285 7868
rect 6144 7828 6150 7840
rect 6273 7837 6285 7840
rect 6319 7837 6331 7871
rect 6273 7831 6331 7837
rect 9122 7828 9128 7880
rect 9180 7868 9186 7880
rect 9401 7871 9459 7877
rect 9401 7868 9413 7871
rect 9180 7840 9413 7868
rect 9180 7828 9186 7840
rect 9401 7837 9413 7840
rect 9447 7837 9459 7871
rect 9401 7831 9459 7837
rect 9582 7828 9588 7880
rect 9640 7828 9646 7880
rect 12526 7828 12532 7880
rect 12584 7828 12590 7880
rect 12636 7877 12664 7908
rect 16853 7905 16865 7939
rect 16899 7936 16911 7939
rect 17678 7936 17684 7948
rect 16899 7908 17684 7936
rect 16899 7905 16911 7908
rect 16853 7899 16911 7905
rect 17678 7896 17684 7908
rect 17736 7896 17742 7948
rect 17880 7908 18368 7936
rect 12621 7871 12679 7877
rect 12621 7837 12633 7871
rect 12667 7837 12679 7871
rect 12621 7831 12679 7837
rect 12710 7828 12716 7880
rect 12768 7828 12774 7880
rect 12894 7828 12900 7880
rect 12952 7828 12958 7880
rect 12986 7828 12992 7880
rect 13044 7828 13050 7880
rect 13814 7828 13820 7880
rect 13872 7868 13878 7880
rect 15746 7868 15752 7880
rect 13872 7840 15752 7868
rect 13872 7828 13878 7840
rect 15746 7828 15752 7840
rect 15804 7828 15810 7880
rect 15930 7828 15936 7880
rect 15988 7877 15994 7880
rect 15988 7871 16037 7877
rect 15988 7837 15991 7871
rect 16025 7837 16037 7871
rect 15988 7831 16037 7837
rect 16117 7871 16175 7877
rect 16117 7837 16129 7871
rect 16163 7868 16175 7871
rect 16942 7868 16948 7880
rect 16163 7840 16948 7868
rect 16163 7837 16175 7840
rect 16117 7831 16175 7837
rect 15988 7828 15994 7831
rect 16942 7828 16948 7840
rect 17000 7828 17006 7880
rect 17034 7828 17040 7880
rect 17092 7828 17098 7880
rect 17126 7828 17132 7880
rect 17184 7868 17190 7880
rect 17497 7871 17555 7877
rect 17497 7868 17509 7871
rect 17184 7840 17509 7868
rect 17184 7828 17190 7840
rect 17497 7837 17509 7840
rect 17543 7837 17555 7871
rect 17497 7831 17555 7837
rect 17586 7828 17592 7880
rect 17644 7828 17650 7880
rect 17770 7828 17776 7880
rect 17828 7828 17834 7880
rect 17880 7877 17908 7908
rect 18156 7877 18276 7878
rect 18340 7877 18368 7908
rect 17865 7871 17923 7877
rect 17865 7837 17877 7871
rect 17911 7837 17923 7871
rect 17865 7831 17923 7837
rect 18141 7871 18276 7877
rect 18141 7837 18153 7871
rect 18187 7850 18276 7871
rect 18187 7837 18199 7850
rect 18141 7831 18199 7837
rect 12253 7803 12311 7809
rect 4479 7772 5764 7800
rect 11822 7772 12204 7800
rect 4479 7769 4491 7772
rect 4433 7763 4491 7769
rect 9493 7735 9551 7741
rect 9493 7701 9505 7735
rect 9539 7732 9551 7735
rect 9950 7732 9956 7744
rect 9539 7704 9956 7732
rect 9539 7701 9551 7704
rect 9493 7695 9551 7701
rect 9950 7692 9956 7704
rect 10008 7732 10014 7744
rect 10594 7732 10600 7744
rect 10008 7704 10600 7732
rect 10008 7692 10014 7704
rect 10594 7692 10600 7704
rect 10652 7692 10658 7744
rect 12176 7732 12204 7772
rect 12253 7769 12265 7803
rect 12299 7800 12311 7803
rect 12342 7800 12348 7812
rect 12299 7772 12348 7800
rect 12299 7769 12311 7772
rect 12253 7763 12311 7769
rect 12342 7760 12348 7772
rect 12400 7760 12406 7812
rect 13722 7760 13728 7812
rect 13780 7760 13786 7812
rect 14182 7800 14188 7812
rect 13832 7772 14188 7800
rect 13170 7732 13176 7744
rect 12176 7704 13176 7732
rect 13170 7692 13176 7704
rect 13228 7692 13234 7744
rect 13354 7692 13360 7744
rect 13412 7692 13418 7744
rect 13525 7735 13583 7741
rect 13525 7701 13537 7735
rect 13571 7732 13583 7735
rect 13832 7732 13860 7772
rect 14182 7760 14188 7772
rect 14240 7760 14246 7812
rect 16574 7760 16580 7812
rect 16632 7800 16638 7812
rect 16761 7803 16819 7809
rect 16761 7800 16773 7803
rect 16632 7772 16773 7800
rect 16632 7760 16638 7772
rect 16761 7769 16773 7772
rect 16807 7769 16819 7803
rect 17880 7800 17908 7831
rect 18248 7812 18276 7850
rect 18325 7871 18383 7877
rect 18325 7837 18337 7871
rect 18371 7837 18383 7871
rect 18325 7831 18383 7837
rect 18414 7828 18420 7880
rect 18472 7828 18478 7880
rect 18506 7828 18512 7880
rect 18564 7828 18570 7880
rect 18598 7828 18604 7880
rect 18656 7828 18662 7880
rect 18782 7828 18788 7880
rect 18840 7828 18846 7880
rect 18874 7828 18880 7880
rect 18932 7828 18938 7880
rect 18046 7800 18052 7812
rect 17880 7772 18052 7800
rect 16761 7763 16819 7769
rect 18046 7760 18052 7772
rect 18104 7760 18110 7812
rect 18230 7760 18236 7812
rect 18288 7800 18294 7812
rect 19150 7800 19156 7812
rect 18288 7772 19156 7800
rect 18288 7760 18294 7772
rect 19150 7760 19156 7772
rect 19208 7760 19214 7812
rect 13571 7704 13860 7732
rect 13571 7701 13583 7704
rect 13525 7695 13583 7701
rect 14550 7692 14556 7744
rect 14608 7732 14614 7744
rect 15194 7732 15200 7744
rect 14608 7704 15200 7732
rect 14608 7692 14614 7704
rect 15194 7692 15200 7704
rect 15252 7692 15258 7744
rect 15930 7692 15936 7744
rect 15988 7732 15994 7744
rect 16666 7732 16672 7744
rect 15988 7704 16672 7732
rect 15988 7692 15994 7704
rect 16666 7692 16672 7704
rect 16724 7692 16730 7744
rect 17034 7692 17040 7744
rect 17092 7732 17098 7744
rect 17313 7735 17371 7741
rect 17313 7732 17325 7735
rect 17092 7704 17325 7732
rect 17092 7692 17098 7704
rect 17313 7701 17325 7704
rect 17359 7701 17371 7735
rect 17313 7695 17371 7701
rect 17402 7692 17408 7744
rect 17460 7732 17466 7744
rect 17957 7735 18015 7741
rect 17957 7732 17969 7735
rect 17460 7704 17969 7732
rect 17460 7692 17466 7704
rect 17957 7701 17969 7704
rect 18003 7701 18015 7735
rect 17957 7695 18015 7701
rect 19058 7692 19064 7744
rect 19116 7692 19122 7744
rect 19242 7692 19248 7744
rect 19300 7692 19306 7744
rect 19352 7732 19380 7976
rect 21192 7948 21220 8035
rect 22186 8032 22192 8084
rect 22244 8072 22250 8084
rect 22244 8044 23520 8072
rect 22244 8032 22250 8044
rect 21266 7964 21272 8016
rect 21324 8004 21330 8016
rect 21545 8007 21603 8013
rect 21545 8004 21557 8007
rect 21324 7976 21557 8004
rect 21324 7964 21330 7976
rect 21545 7973 21557 7976
rect 21591 7973 21603 8007
rect 23382 8004 23388 8016
rect 21545 7967 21603 7973
rect 22940 7976 23388 8004
rect 19702 7896 19708 7948
rect 19760 7936 19766 7948
rect 20809 7939 20867 7945
rect 20809 7936 20821 7939
rect 19760 7908 20821 7936
rect 19760 7896 19766 7908
rect 20809 7905 20821 7908
rect 20855 7905 20867 7939
rect 20809 7899 20867 7905
rect 21174 7896 21180 7948
rect 21232 7896 21238 7948
rect 21560 7936 21588 7967
rect 21560 7908 22048 7936
rect 19518 7828 19524 7880
rect 19576 7828 19582 7880
rect 19610 7828 19616 7880
rect 19668 7868 19674 7880
rect 19797 7871 19855 7877
rect 19797 7868 19809 7871
rect 19668 7840 19809 7868
rect 19668 7828 19674 7840
rect 19797 7837 19809 7840
rect 19843 7837 19855 7871
rect 19797 7831 19855 7837
rect 19978 7828 19984 7880
rect 20036 7828 20042 7880
rect 20257 7871 20315 7877
rect 20257 7837 20269 7871
rect 20303 7837 20315 7871
rect 20257 7831 20315 7837
rect 20349 7871 20407 7877
rect 20349 7837 20361 7871
rect 20395 7868 20407 7871
rect 20438 7868 20444 7880
rect 20395 7840 20444 7868
rect 20395 7837 20407 7840
rect 20349 7831 20407 7837
rect 19426 7760 19432 7812
rect 19484 7800 19490 7812
rect 19996 7800 20024 7828
rect 19484 7772 20024 7800
rect 20272 7800 20300 7831
rect 20438 7828 20444 7840
rect 20496 7828 20502 7880
rect 20530 7828 20536 7880
rect 20588 7828 20594 7880
rect 20622 7828 20628 7880
rect 20680 7828 20686 7880
rect 20901 7871 20959 7877
rect 20901 7837 20913 7871
rect 20947 7868 20959 7871
rect 21082 7868 21088 7880
rect 20947 7840 21088 7868
rect 20947 7837 20959 7840
rect 20901 7831 20959 7837
rect 21082 7828 21088 7840
rect 21140 7868 21146 7880
rect 21542 7868 21548 7880
rect 21140 7840 21548 7868
rect 21140 7828 21146 7840
rect 21542 7828 21548 7840
rect 21600 7828 21606 7880
rect 22020 7877 22048 7908
rect 22940 7877 22968 7976
rect 23382 7964 23388 7976
rect 23440 7964 23446 8016
rect 23492 8004 23520 8044
rect 23750 8032 23756 8084
rect 23808 8032 23814 8084
rect 24857 8075 24915 8081
rect 24857 8041 24869 8075
rect 24903 8072 24915 8075
rect 25038 8072 25044 8084
rect 24903 8044 25044 8072
rect 24903 8041 24915 8044
rect 24857 8035 24915 8041
rect 25038 8032 25044 8044
rect 25096 8032 25102 8084
rect 23842 8004 23848 8016
rect 23492 7976 23848 8004
rect 23842 7964 23848 7976
rect 23900 7964 23906 8016
rect 24302 7964 24308 8016
rect 24360 8004 24366 8016
rect 24397 8007 24455 8013
rect 24397 8004 24409 8007
rect 24360 7976 24409 8004
rect 24360 7964 24366 7976
rect 24397 7973 24409 7976
rect 24443 7973 24455 8007
rect 24397 7967 24455 7973
rect 23293 7939 23351 7945
rect 23293 7905 23305 7939
rect 23339 7936 23351 7939
rect 23474 7936 23480 7948
rect 23339 7908 23480 7936
rect 23339 7905 23351 7908
rect 23293 7899 23351 7905
rect 23474 7896 23480 7908
rect 23532 7896 23538 7948
rect 24762 7936 24768 7948
rect 23676 7908 24768 7936
rect 22005 7871 22063 7877
rect 22005 7837 22017 7871
rect 22051 7837 22063 7871
rect 22005 7831 22063 7837
rect 22925 7871 22983 7877
rect 22925 7837 22937 7871
rect 22971 7837 22983 7871
rect 22925 7831 22983 7837
rect 23109 7871 23167 7877
rect 23109 7837 23121 7871
rect 23155 7868 23167 7871
rect 23385 7871 23443 7877
rect 23385 7868 23397 7871
rect 23155 7840 23397 7868
rect 23155 7837 23167 7840
rect 23109 7831 23167 7837
rect 23385 7837 23397 7840
rect 23431 7868 23443 7871
rect 23676 7868 23704 7908
rect 24762 7896 24768 7908
rect 24820 7896 24826 7948
rect 23431 7840 23704 7868
rect 23431 7837 23443 7840
rect 23385 7831 23443 7837
rect 23750 7828 23756 7880
rect 23808 7868 23814 7880
rect 24029 7871 24087 7877
rect 24029 7868 24041 7871
rect 23808 7840 24041 7868
rect 23808 7828 23814 7840
rect 24029 7837 24041 7840
rect 24075 7837 24087 7871
rect 24029 7831 24087 7837
rect 24118 7828 24124 7880
rect 24176 7828 24182 7880
rect 25041 7871 25099 7877
rect 25041 7837 25053 7871
rect 25087 7868 25099 7871
rect 25682 7868 25688 7880
rect 25087 7840 25688 7868
rect 25087 7837 25099 7840
rect 25041 7831 25099 7837
rect 25682 7828 25688 7840
rect 25740 7868 25746 7880
rect 27706 7868 27712 7880
rect 25740 7840 27712 7868
rect 25740 7828 25746 7840
rect 27706 7828 27712 7840
rect 27764 7828 27770 7880
rect 21634 7800 21640 7812
rect 20272 7772 21640 7800
rect 19484 7760 19490 7772
rect 21634 7760 21640 7772
rect 21692 7760 21698 7812
rect 21821 7803 21879 7809
rect 21821 7769 21833 7803
rect 21867 7800 21879 7803
rect 23290 7800 23296 7812
rect 21867 7772 23296 7800
rect 21867 7769 21879 7772
rect 21821 7763 21879 7769
rect 23290 7760 23296 7772
rect 23348 7760 23354 7812
rect 24581 7803 24639 7809
rect 24581 7769 24593 7803
rect 24627 7800 24639 7803
rect 27614 7800 27620 7812
rect 24627 7772 27620 7800
rect 24627 7769 24639 7772
rect 24581 7763 24639 7769
rect 27614 7760 27620 7772
rect 27672 7760 27678 7812
rect 21726 7732 21732 7744
rect 19352 7704 21732 7732
rect 21726 7692 21732 7704
rect 21784 7692 21790 7744
rect 22738 7692 22744 7744
rect 22796 7692 22802 7744
rect 23750 7692 23756 7744
rect 23808 7732 23814 7744
rect 23845 7735 23903 7741
rect 23845 7732 23857 7735
rect 23808 7704 23857 7732
rect 23808 7692 23814 7704
rect 23845 7701 23857 7704
rect 23891 7701 23903 7735
rect 23845 7695 23903 7701
rect 1104 7642 28152 7664
rect 1104 7590 4874 7642
rect 4926 7590 4938 7642
rect 4990 7590 5002 7642
rect 5054 7590 5066 7642
rect 5118 7590 5130 7642
rect 5182 7590 28152 7642
rect 1104 7568 28152 7590
rect 4709 7531 4767 7537
rect 4709 7497 4721 7531
rect 4755 7528 4767 7531
rect 4798 7528 4804 7540
rect 4755 7500 4804 7528
rect 4755 7497 4767 7500
rect 4709 7491 4767 7497
rect 4798 7488 4804 7500
rect 4856 7488 4862 7540
rect 5258 7488 5264 7540
rect 5316 7488 5322 7540
rect 7929 7531 7987 7537
rect 7929 7497 7941 7531
rect 7975 7528 7987 7531
rect 8018 7528 8024 7540
rect 7975 7500 8024 7528
rect 7975 7497 7987 7500
rect 7929 7491 7987 7497
rect 8018 7488 8024 7500
rect 8076 7488 8082 7540
rect 8294 7488 8300 7540
rect 8352 7528 8358 7540
rect 8846 7528 8852 7540
rect 8352 7500 8852 7528
rect 8352 7488 8358 7500
rect 8846 7488 8852 7500
rect 8904 7488 8910 7540
rect 9766 7528 9772 7540
rect 9324 7500 9772 7528
rect 5276 7460 5304 7488
rect 4632 7432 5304 7460
rect 6472 7432 7696 7460
rect 4632 7401 4660 7432
rect 4617 7395 4675 7401
rect 4617 7361 4629 7395
rect 4663 7361 4675 7395
rect 4617 7355 4675 7361
rect 4801 7395 4859 7401
rect 4801 7361 4813 7395
rect 4847 7392 4859 7395
rect 5261 7395 5319 7401
rect 4847 7364 4936 7392
rect 4847 7361 4859 7364
rect 4801 7355 4859 7361
rect 4908 7197 4936 7364
rect 5261 7361 5273 7395
rect 5307 7392 5319 7395
rect 5534 7392 5540 7404
rect 5307 7364 5540 7392
rect 5307 7361 5319 7364
rect 5261 7355 5319 7361
rect 5534 7352 5540 7364
rect 5592 7352 5598 7404
rect 5721 7395 5779 7401
rect 5721 7361 5733 7395
rect 5767 7361 5779 7395
rect 5721 7355 5779 7361
rect 5353 7327 5411 7333
rect 5353 7293 5365 7327
rect 5399 7293 5411 7327
rect 5353 7287 5411 7293
rect 5368 7256 5396 7287
rect 5442 7284 5448 7336
rect 5500 7324 5506 7336
rect 5629 7327 5687 7333
rect 5629 7324 5641 7327
rect 5500 7296 5641 7324
rect 5500 7284 5506 7296
rect 5629 7293 5641 7296
rect 5675 7293 5687 7327
rect 5736 7324 5764 7355
rect 5810 7352 5816 7404
rect 5868 7392 5874 7404
rect 6365 7395 6423 7401
rect 6365 7392 6377 7395
rect 5868 7364 6377 7392
rect 5868 7352 5874 7364
rect 6365 7361 6377 7364
rect 6411 7392 6423 7395
rect 6472 7392 6500 7432
rect 6411 7364 6500 7392
rect 6411 7361 6423 7364
rect 6365 7355 6423 7361
rect 6546 7352 6552 7404
rect 6604 7352 6610 7404
rect 6457 7327 6515 7333
rect 6457 7324 6469 7327
rect 5736 7296 6469 7324
rect 5629 7287 5687 7293
rect 6457 7293 6469 7296
rect 6503 7293 6515 7327
rect 6457 7287 6515 7293
rect 6089 7259 6147 7265
rect 5368 7228 5672 7256
rect 4893 7191 4951 7197
rect 4893 7157 4905 7191
rect 4939 7188 4951 7191
rect 5534 7188 5540 7200
rect 4939 7160 5540 7188
rect 4939 7157 4951 7160
rect 4893 7151 4951 7157
rect 5534 7148 5540 7160
rect 5592 7148 5598 7200
rect 5644 7188 5672 7228
rect 6089 7225 6101 7259
rect 6135 7256 6147 7259
rect 7558 7256 7564 7268
rect 6135 7228 7564 7256
rect 6135 7225 6147 7228
rect 6089 7219 6147 7225
rect 7558 7216 7564 7228
rect 7616 7216 7622 7268
rect 7668 7256 7696 7432
rect 8018 7352 8024 7404
rect 8076 7392 8082 7404
rect 8113 7395 8171 7401
rect 8113 7392 8125 7395
rect 8076 7364 8125 7392
rect 8076 7352 8082 7364
rect 8113 7361 8125 7364
rect 8159 7361 8171 7395
rect 8113 7355 8171 7361
rect 8386 7352 8392 7404
rect 8444 7352 8450 7404
rect 8478 7352 8484 7404
rect 8536 7352 8542 7404
rect 8570 7352 8576 7404
rect 8628 7392 8634 7404
rect 8665 7395 8723 7401
rect 8665 7392 8677 7395
rect 8628 7364 8677 7392
rect 8628 7352 8634 7364
rect 8665 7361 8677 7364
rect 8711 7392 8723 7395
rect 9030 7392 9036 7404
rect 8711 7364 9036 7392
rect 8711 7361 8723 7364
rect 8665 7355 8723 7361
rect 9030 7352 9036 7364
rect 9088 7352 9094 7404
rect 9122 7352 9128 7404
rect 9180 7352 9186 7404
rect 9217 7395 9275 7401
rect 9217 7361 9229 7395
rect 9263 7361 9275 7395
rect 9324 7392 9352 7500
rect 9766 7488 9772 7500
rect 9824 7488 9830 7540
rect 12158 7488 12164 7540
rect 12216 7488 12222 7540
rect 12713 7531 12771 7537
rect 12713 7497 12725 7531
rect 12759 7528 12771 7531
rect 12986 7528 12992 7540
rect 12759 7500 12992 7528
rect 12759 7497 12771 7500
rect 12713 7491 12771 7497
rect 12986 7488 12992 7500
rect 13044 7488 13050 7540
rect 14090 7488 14096 7540
rect 14148 7488 14154 7540
rect 14550 7488 14556 7540
rect 14608 7488 14614 7540
rect 14921 7531 14979 7537
rect 14921 7497 14933 7531
rect 14967 7528 14979 7531
rect 15010 7528 15016 7540
rect 14967 7500 15016 7528
rect 14967 7497 14979 7500
rect 14921 7491 14979 7497
rect 15010 7488 15016 7500
rect 15068 7488 15074 7540
rect 16206 7488 16212 7540
rect 16264 7488 16270 7540
rect 17678 7488 17684 7540
rect 17736 7528 17742 7540
rect 17865 7531 17923 7537
rect 17865 7528 17877 7531
rect 17736 7500 17877 7528
rect 17736 7488 17742 7500
rect 17865 7497 17877 7500
rect 17911 7497 17923 7531
rect 17865 7491 17923 7497
rect 18046 7488 18052 7540
rect 18104 7488 18110 7540
rect 18138 7488 18144 7540
rect 18196 7528 18202 7540
rect 18325 7531 18383 7537
rect 18325 7528 18337 7531
rect 18196 7500 18337 7528
rect 18196 7488 18202 7500
rect 18325 7497 18337 7500
rect 18371 7497 18383 7531
rect 18325 7491 18383 7497
rect 18414 7488 18420 7540
rect 18472 7528 18478 7540
rect 20070 7528 20076 7540
rect 18472 7500 20076 7528
rect 18472 7488 18478 7500
rect 20070 7488 20076 7500
rect 20128 7488 20134 7540
rect 20530 7488 20536 7540
rect 20588 7528 20594 7540
rect 20625 7531 20683 7537
rect 20625 7528 20637 7531
rect 20588 7500 20637 7528
rect 20588 7488 20594 7500
rect 20625 7497 20637 7500
rect 20671 7497 20683 7531
rect 22557 7531 22615 7537
rect 22557 7528 22569 7531
rect 20625 7491 20683 7497
rect 20824 7500 22569 7528
rect 9401 7463 9459 7469
rect 9401 7429 9413 7463
rect 9447 7460 9459 7463
rect 10413 7463 10471 7469
rect 10413 7460 10425 7463
rect 9447 7432 10425 7460
rect 9447 7429 9459 7432
rect 9401 7423 9459 7429
rect 10413 7429 10425 7432
rect 10459 7429 10471 7463
rect 10413 7423 10471 7429
rect 10594 7420 10600 7472
rect 10652 7420 10658 7472
rect 10781 7463 10839 7469
rect 10781 7429 10793 7463
rect 10827 7460 10839 7463
rect 10870 7460 10876 7472
rect 10827 7432 10876 7460
rect 10827 7429 10839 7432
rect 10781 7423 10839 7429
rect 10870 7420 10876 7432
rect 10928 7420 10934 7472
rect 11517 7463 11575 7469
rect 11517 7429 11529 7463
rect 11563 7460 11575 7463
rect 12434 7460 12440 7472
rect 11563 7432 12440 7460
rect 11563 7429 11575 7432
rect 11517 7423 11575 7429
rect 12434 7420 12440 7432
rect 12492 7420 12498 7472
rect 13078 7460 13084 7472
rect 13004 7432 13084 7460
rect 9493 7395 9551 7401
rect 9493 7392 9505 7395
rect 9324 7364 9505 7392
rect 9217 7355 9275 7361
rect 9493 7361 9505 7364
rect 9539 7361 9551 7395
rect 9493 7355 9551 7361
rect 9232 7324 9260 7355
rect 9674 7352 9680 7404
rect 9732 7352 9738 7404
rect 9861 7395 9919 7401
rect 9861 7361 9873 7395
rect 9907 7392 9919 7395
rect 9953 7395 10011 7401
rect 9953 7392 9965 7395
rect 9907 7364 9965 7392
rect 9907 7361 9919 7364
rect 9861 7355 9919 7361
rect 9953 7361 9965 7364
rect 9999 7361 10011 7395
rect 9953 7355 10011 7361
rect 10137 7395 10195 7401
rect 10137 7361 10149 7395
rect 10183 7361 10195 7395
rect 10137 7355 10195 7361
rect 10321 7395 10379 7401
rect 10321 7361 10333 7395
rect 10367 7392 10379 7395
rect 10686 7392 10692 7404
rect 10367 7364 10692 7392
rect 10367 7361 10379 7364
rect 10321 7355 10379 7361
rect 9582 7324 9588 7336
rect 9232 7296 9588 7324
rect 9582 7284 9588 7296
rect 9640 7324 9646 7336
rect 10152 7324 10180 7355
rect 10686 7352 10692 7364
rect 10744 7352 10750 7404
rect 11606 7352 11612 7404
rect 11664 7352 11670 7404
rect 11882 7352 11888 7404
rect 11940 7352 11946 7404
rect 13004 7401 13032 7432
rect 13078 7420 13084 7432
rect 13136 7460 13142 7472
rect 13136 7432 14688 7460
rect 13136 7420 13142 7432
rect 12989 7395 13047 7401
rect 12989 7361 13001 7395
rect 13035 7361 13047 7395
rect 12989 7355 13047 7361
rect 13173 7395 13231 7401
rect 13173 7361 13185 7395
rect 13219 7392 13231 7395
rect 13354 7392 13360 7404
rect 13219 7364 13360 7392
rect 13219 7361 13231 7364
rect 13173 7355 13231 7361
rect 13354 7352 13360 7364
rect 13412 7352 13418 7404
rect 13446 7352 13452 7404
rect 13504 7352 13510 7404
rect 13541 7395 13599 7401
rect 13541 7361 13553 7395
rect 13587 7361 13599 7395
rect 13541 7355 13599 7361
rect 9640 7296 10180 7324
rect 9640 7284 9646 7296
rect 11624 7256 11652 7352
rect 11698 7284 11704 7336
rect 11756 7324 11762 7336
rect 11977 7327 12035 7333
rect 11977 7324 11989 7327
rect 11756 7296 11989 7324
rect 11756 7284 11762 7296
rect 11977 7293 11989 7296
rect 12023 7324 12035 7327
rect 13556 7324 13584 7355
rect 13814 7352 13820 7404
rect 13872 7352 13878 7404
rect 13906 7352 13912 7404
rect 13964 7352 13970 7404
rect 14461 7395 14519 7401
rect 14461 7361 14473 7395
rect 14507 7392 14519 7395
rect 14550 7392 14556 7404
rect 14507 7364 14556 7392
rect 14507 7361 14519 7364
rect 14461 7355 14519 7361
rect 14550 7352 14556 7364
rect 14608 7352 14614 7404
rect 12023 7296 13584 7324
rect 13633 7327 13691 7333
rect 12023 7293 12035 7296
rect 11977 7287 12035 7293
rect 13633 7293 13645 7327
rect 13679 7324 13691 7327
rect 13722 7324 13728 7336
rect 13679 7296 13728 7324
rect 13679 7293 13691 7296
rect 13633 7287 13691 7293
rect 13722 7284 13728 7296
rect 13780 7284 13786 7336
rect 14660 7333 14688 7432
rect 14734 7420 14740 7472
rect 14792 7460 14798 7472
rect 14792 7432 14964 7460
rect 14792 7420 14798 7432
rect 14826 7352 14832 7404
rect 14884 7352 14890 7404
rect 14936 7392 14964 7432
rect 15194 7420 15200 7472
rect 15252 7460 15258 7472
rect 15657 7463 15715 7469
rect 15657 7460 15669 7463
rect 15252 7432 15669 7460
rect 15252 7420 15258 7432
rect 15657 7429 15669 7432
rect 15703 7429 15715 7463
rect 16224 7460 16252 7488
rect 18432 7460 18460 7488
rect 15657 7423 15715 7429
rect 16132 7432 16252 7460
rect 17512 7432 18460 7460
rect 15102 7392 15108 7404
rect 14936 7364 15108 7392
rect 15102 7352 15108 7364
rect 15160 7352 15166 7404
rect 15289 7395 15347 7401
rect 15289 7361 15301 7395
rect 15335 7361 15347 7395
rect 15289 7355 15347 7361
rect 14645 7327 14703 7333
rect 14645 7293 14657 7327
rect 14691 7324 14703 7327
rect 15304 7324 15332 7355
rect 15378 7352 15384 7404
rect 15436 7392 15442 7404
rect 15473 7395 15531 7401
rect 15473 7392 15485 7395
rect 15436 7364 15485 7392
rect 15436 7352 15442 7364
rect 15473 7361 15485 7364
rect 15519 7361 15531 7395
rect 15473 7355 15531 7361
rect 15562 7352 15568 7404
rect 15620 7352 15626 7404
rect 15838 7352 15844 7404
rect 15896 7352 15902 7404
rect 15930 7352 15936 7404
rect 15988 7352 15994 7404
rect 16132 7401 16160 7432
rect 16117 7395 16175 7401
rect 16117 7361 16129 7395
rect 16163 7361 16175 7395
rect 16117 7355 16175 7361
rect 16206 7352 16212 7404
rect 16264 7352 16270 7404
rect 16301 7395 16359 7401
rect 16301 7361 16313 7395
rect 16347 7392 16359 7395
rect 16574 7392 16580 7404
rect 16347 7364 16580 7392
rect 16347 7361 16359 7364
rect 16301 7355 16359 7361
rect 16574 7352 16580 7364
rect 16632 7352 16638 7404
rect 16758 7352 16764 7404
rect 16816 7352 16822 7404
rect 16853 7395 16911 7401
rect 16853 7361 16865 7395
rect 16899 7392 16911 7395
rect 17034 7392 17040 7404
rect 16899 7364 17040 7392
rect 16899 7361 16911 7364
rect 16853 7355 16911 7361
rect 17034 7352 17040 7364
rect 17092 7352 17098 7404
rect 17129 7395 17187 7401
rect 17129 7361 17141 7395
rect 17175 7392 17187 7395
rect 17402 7392 17408 7404
rect 17175 7364 17408 7392
rect 17175 7361 17187 7364
rect 17129 7355 17187 7361
rect 17402 7352 17408 7364
rect 17460 7352 17466 7404
rect 14691 7296 15332 7324
rect 16224 7324 16252 7352
rect 16393 7327 16451 7333
rect 16393 7324 16405 7327
rect 16224 7296 16405 7324
rect 14691 7293 14703 7296
rect 14645 7287 14703 7293
rect 14366 7256 14372 7268
rect 7668 7228 11652 7256
rect 11716 7228 14372 7256
rect 6546 7188 6552 7200
rect 5644 7160 6552 7188
rect 6546 7148 6552 7160
rect 6604 7148 6610 7200
rect 9030 7148 9036 7200
rect 9088 7188 9094 7200
rect 11716 7188 11744 7228
rect 14366 7216 14372 7228
rect 14424 7216 14430 7268
rect 15304 7256 15332 7296
rect 16393 7293 16405 7296
rect 16439 7293 16451 7327
rect 16393 7287 16451 7293
rect 16945 7327 17003 7333
rect 16945 7293 16957 7327
rect 16991 7293 17003 7327
rect 16945 7287 17003 7293
rect 17221 7327 17279 7333
rect 17221 7293 17233 7327
rect 17267 7293 17279 7327
rect 17221 7287 17279 7293
rect 16850 7256 16856 7268
rect 15304 7228 16856 7256
rect 16850 7216 16856 7228
rect 16908 7256 16914 7268
rect 16960 7256 16988 7287
rect 16908 7228 16988 7256
rect 16908 7216 16914 7228
rect 17034 7216 17040 7268
rect 17092 7256 17098 7268
rect 17129 7259 17187 7265
rect 17129 7256 17141 7259
rect 17092 7228 17141 7256
rect 17092 7216 17098 7228
rect 17129 7225 17141 7228
rect 17175 7256 17187 7259
rect 17236 7256 17264 7287
rect 17310 7284 17316 7336
rect 17368 7284 17374 7336
rect 17175 7228 17264 7256
rect 17175 7225 17187 7228
rect 17129 7219 17187 7225
rect 9088 7160 11744 7188
rect 9088 7148 9094 7160
rect 12434 7148 12440 7200
rect 12492 7188 12498 7200
rect 12986 7188 12992 7200
rect 12492 7160 12992 7188
rect 12492 7148 12498 7160
rect 12986 7148 12992 7160
rect 13044 7148 13050 7200
rect 13078 7148 13084 7200
rect 13136 7148 13142 7200
rect 13262 7148 13268 7200
rect 13320 7148 13326 7200
rect 14829 7191 14887 7197
rect 14829 7157 14841 7191
rect 14875 7188 14887 7191
rect 16022 7188 16028 7200
rect 14875 7160 16028 7188
rect 14875 7157 14887 7160
rect 14829 7151 14887 7157
rect 16022 7148 16028 7160
rect 16080 7148 16086 7200
rect 16298 7148 16304 7200
rect 16356 7188 16362 7200
rect 17512 7188 17540 7432
rect 18506 7420 18512 7472
rect 18564 7460 18570 7472
rect 20088 7460 20116 7488
rect 20257 7463 20315 7469
rect 18564 7432 19564 7460
rect 20088 7432 20208 7460
rect 18564 7420 18570 7432
rect 17586 7352 17592 7404
rect 17644 7352 17650 7404
rect 17681 7395 17739 7401
rect 17681 7361 17693 7395
rect 17727 7392 17739 7395
rect 17862 7392 17868 7404
rect 17727 7364 17868 7392
rect 17727 7361 17739 7364
rect 17681 7355 17739 7361
rect 17862 7352 17868 7364
rect 17920 7352 17926 7404
rect 17954 7352 17960 7404
rect 18012 7392 18018 7404
rect 18141 7395 18199 7401
rect 18141 7392 18153 7395
rect 18012 7364 18153 7392
rect 18012 7352 18018 7364
rect 18141 7361 18153 7364
rect 18187 7361 18199 7395
rect 18141 7355 18199 7361
rect 18156 7324 18184 7355
rect 18230 7352 18236 7404
rect 18288 7352 18294 7404
rect 19058 7352 19064 7404
rect 19116 7352 19122 7404
rect 19536 7401 19564 7432
rect 20180 7401 20208 7432
rect 20257 7429 20269 7463
rect 20303 7460 20315 7463
rect 20824 7460 20852 7500
rect 22557 7497 22569 7500
rect 22603 7497 22615 7531
rect 22557 7491 22615 7497
rect 23290 7488 23296 7540
rect 23348 7488 23354 7540
rect 24762 7488 24768 7540
rect 24820 7528 24826 7540
rect 25225 7531 25283 7537
rect 25225 7528 25237 7531
rect 24820 7500 25237 7528
rect 24820 7488 24826 7500
rect 25225 7497 25237 7500
rect 25271 7497 25283 7531
rect 25225 7491 25283 7497
rect 20303 7432 20852 7460
rect 20303 7429 20315 7432
rect 20257 7423 20315 7429
rect 20732 7401 20760 7432
rect 21174 7420 21180 7472
rect 21232 7460 21238 7472
rect 21232 7432 22232 7460
rect 21232 7420 21238 7432
rect 19521 7395 19579 7401
rect 19521 7361 19533 7395
rect 19567 7361 19579 7395
rect 19521 7355 19579 7361
rect 20165 7395 20223 7401
rect 20165 7361 20177 7395
rect 20211 7361 20223 7395
rect 20165 7355 20223 7361
rect 20441 7395 20499 7401
rect 20441 7361 20453 7395
rect 20487 7361 20499 7395
rect 20441 7355 20499 7361
rect 20717 7395 20775 7401
rect 20717 7361 20729 7395
rect 20763 7361 20775 7395
rect 20717 7355 20775 7361
rect 18598 7324 18604 7336
rect 18156 7296 18604 7324
rect 18598 7284 18604 7296
rect 18656 7284 18662 7336
rect 19242 7284 19248 7336
rect 19300 7284 19306 7336
rect 19705 7327 19763 7333
rect 19705 7293 19717 7327
rect 19751 7293 19763 7327
rect 19705 7287 19763 7293
rect 16356 7160 17540 7188
rect 19720 7188 19748 7287
rect 19794 7284 19800 7336
rect 19852 7324 19858 7336
rect 20456 7324 20484 7355
rect 20806 7352 20812 7404
rect 20864 7352 20870 7404
rect 20898 7352 20904 7404
rect 20956 7392 20962 7404
rect 20993 7395 21051 7401
rect 20993 7392 21005 7395
rect 20956 7364 21005 7392
rect 20956 7352 20962 7364
rect 20993 7361 21005 7364
rect 21039 7361 21051 7395
rect 20993 7355 21051 7361
rect 21082 7352 21088 7404
rect 21140 7352 21146 7404
rect 21361 7395 21419 7401
rect 21361 7361 21373 7395
rect 21407 7361 21419 7395
rect 21545 7395 21603 7401
rect 21545 7392 21557 7395
rect 21361 7355 21419 7361
rect 21468 7364 21557 7392
rect 19852 7296 20484 7324
rect 19852 7284 19858 7296
rect 20530 7284 20536 7336
rect 20588 7324 20594 7336
rect 21376 7324 21404 7355
rect 20588 7296 21404 7324
rect 20588 7284 20594 7296
rect 20438 7216 20444 7268
rect 20496 7256 20502 7268
rect 21269 7259 21327 7265
rect 21269 7256 21281 7259
rect 20496 7228 21281 7256
rect 20496 7216 20502 7228
rect 21269 7225 21281 7228
rect 21315 7256 21327 7259
rect 21468 7256 21496 7364
rect 21545 7361 21557 7364
rect 21591 7361 21603 7395
rect 21545 7355 21603 7361
rect 21634 7352 21640 7404
rect 21692 7392 21698 7404
rect 21821 7395 21879 7401
rect 21821 7392 21833 7395
rect 21692 7364 21833 7392
rect 21692 7352 21698 7364
rect 21821 7361 21833 7364
rect 21867 7361 21879 7395
rect 21821 7355 21879 7361
rect 22002 7352 22008 7404
rect 22060 7352 22066 7404
rect 22204 7401 22232 7432
rect 23750 7420 23756 7472
rect 23808 7420 23814 7472
rect 25038 7460 25044 7472
rect 24978 7432 25044 7460
rect 25038 7420 25044 7432
rect 25096 7420 25102 7472
rect 22189 7395 22247 7401
rect 22189 7361 22201 7395
rect 22235 7361 22247 7395
rect 22189 7355 22247 7361
rect 22278 7352 22284 7404
rect 22336 7352 22342 7404
rect 22462 7352 22468 7404
rect 22520 7352 22526 7404
rect 23382 7352 23388 7404
rect 23440 7352 23446 7404
rect 23474 7352 23480 7404
rect 23532 7352 23538 7404
rect 21726 7284 21732 7336
rect 21784 7324 21790 7336
rect 23400 7324 23428 7352
rect 21784 7296 23428 7324
rect 21784 7284 21790 7296
rect 21315 7228 21496 7256
rect 22097 7259 22155 7265
rect 21315 7225 21327 7228
rect 21269 7219 21327 7225
rect 22097 7225 22109 7259
rect 22143 7256 22155 7259
rect 22370 7256 22376 7268
rect 22143 7228 22376 7256
rect 22143 7225 22155 7228
rect 22097 7219 22155 7225
rect 22370 7216 22376 7228
rect 22428 7216 22434 7268
rect 21174 7188 21180 7200
rect 19720 7160 21180 7188
rect 16356 7148 16362 7160
rect 21174 7148 21180 7160
rect 21232 7148 21238 7200
rect 21358 7148 21364 7200
rect 21416 7148 21422 7200
rect 1104 7098 28152 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 28152 7098
rect 1104 7024 28152 7046
rect 8018 6944 8024 6996
rect 8076 6944 8082 6996
rect 9122 6944 9128 6996
rect 9180 6984 9186 6996
rect 9401 6987 9459 6993
rect 9401 6984 9413 6987
rect 9180 6956 9413 6984
rect 9180 6944 9186 6956
rect 9401 6953 9413 6956
rect 9447 6953 9459 6987
rect 9401 6947 9459 6953
rect 9582 6944 9588 6996
rect 9640 6984 9646 6996
rect 9677 6987 9735 6993
rect 9677 6984 9689 6987
rect 9640 6956 9689 6984
rect 9640 6944 9646 6956
rect 9677 6953 9689 6956
rect 9723 6953 9735 6987
rect 12437 6987 12495 6993
rect 12437 6984 12449 6987
rect 9677 6947 9735 6953
rect 12176 6956 12449 6984
rect 5258 6876 5264 6928
rect 5316 6916 5322 6928
rect 5316 6888 5672 6916
rect 5316 6876 5322 6888
rect 5534 6808 5540 6860
rect 5592 6808 5598 6860
rect 5644 6789 5672 6888
rect 7558 6876 7564 6928
rect 7616 6916 7622 6928
rect 8113 6919 8171 6925
rect 8113 6916 8125 6919
rect 7616 6888 8125 6916
rect 7616 6876 7622 6888
rect 8113 6885 8125 6888
rect 8159 6885 8171 6919
rect 8113 6879 8171 6885
rect 8478 6876 8484 6928
rect 8536 6916 8542 6928
rect 8536 6888 9628 6916
rect 8536 6876 8542 6888
rect 7653 6851 7711 6857
rect 7653 6817 7665 6851
rect 7699 6817 7711 6851
rect 7653 6811 7711 6817
rect 5629 6783 5687 6789
rect 5629 6749 5641 6783
rect 5675 6749 5687 6783
rect 5629 6743 5687 6749
rect 7558 6740 7564 6792
rect 7616 6740 7622 6792
rect 7668 6712 7696 6811
rect 8386 6808 8392 6860
rect 8444 6848 8450 6860
rect 9033 6851 9091 6857
rect 9033 6848 9045 6851
rect 8444 6820 9045 6848
rect 8444 6808 8450 6820
rect 9033 6817 9045 6820
rect 9079 6817 9091 6851
rect 9600 6848 9628 6888
rect 11882 6876 11888 6928
rect 11940 6876 11946 6928
rect 12176 6848 12204 6956
rect 12437 6953 12449 6956
rect 12483 6984 12495 6987
rect 12894 6984 12900 6996
rect 12483 6956 12900 6984
rect 12483 6953 12495 6956
rect 12437 6947 12495 6953
rect 12894 6944 12900 6956
rect 12952 6944 12958 6996
rect 13078 6944 13084 6996
rect 13136 6984 13142 6996
rect 13633 6987 13691 6993
rect 13633 6984 13645 6987
rect 13136 6956 13645 6984
rect 13136 6944 13142 6956
rect 13633 6953 13645 6956
rect 13679 6953 13691 6987
rect 13633 6947 13691 6953
rect 15010 6944 15016 6996
rect 15068 6944 15074 6996
rect 15102 6944 15108 6996
rect 15160 6984 15166 6996
rect 15197 6987 15255 6993
rect 15197 6984 15209 6987
rect 15160 6956 15209 6984
rect 15160 6944 15166 6956
rect 15197 6953 15209 6956
rect 15243 6953 15255 6987
rect 15197 6947 15255 6953
rect 15289 6987 15347 6993
rect 15289 6953 15301 6987
rect 15335 6984 15347 6987
rect 15378 6984 15384 6996
rect 15335 6956 15384 6984
rect 15335 6953 15347 6956
rect 15289 6947 15347 6953
rect 15378 6944 15384 6956
rect 15436 6944 15442 6996
rect 15746 6944 15752 6996
rect 15804 6984 15810 6996
rect 15933 6987 15991 6993
rect 15933 6984 15945 6987
rect 15804 6956 15945 6984
rect 15804 6944 15810 6956
rect 15933 6953 15945 6956
rect 15979 6953 15991 6987
rect 15933 6947 15991 6953
rect 16666 6944 16672 6996
rect 16724 6984 16730 6996
rect 17310 6984 17316 6996
rect 16724 6956 17316 6984
rect 16724 6944 16730 6956
rect 17310 6944 17316 6956
rect 17368 6944 17374 6996
rect 17586 6944 17592 6996
rect 17644 6984 17650 6996
rect 20330 6987 20388 6993
rect 20330 6984 20342 6987
rect 17644 6956 20342 6984
rect 17644 6944 17650 6956
rect 20330 6953 20342 6956
rect 20376 6984 20388 6987
rect 21358 6984 21364 6996
rect 20376 6956 21364 6984
rect 20376 6953 20388 6956
rect 20330 6947 20388 6953
rect 21358 6944 21364 6956
rect 21416 6944 21422 6996
rect 21542 6944 21548 6996
rect 21600 6984 21606 6996
rect 21821 6987 21879 6993
rect 21821 6984 21833 6987
rect 21600 6956 21833 6984
rect 21600 6944 21606 6956
rect 21821 6953 21833 6956
rect 21867 6984 21879 6987
rect 22462 6984 22468 6996
rect 21867 6956 22468 6984
rect 21867 6953 21879 6956
rect 21821 6947 21879 6953
rect 22462 6944 22468 6956
rect 22520 6944 22526 6996
rect 12250 6876 12256 6928
rect 12308 6916 12314 6928
rect 12308 6888 12572 6916
rect 12308 6876 12314 6888
rect 9600 6820 10180 6848
rect 9033 6811 9091 6817
rect 8570 6740 8576 6792
rect 8628 6740 8634 6792
rect 8754 6740 8760 6792
rect 8812 6740 8818 6792
rect 8846 6740 8852 6792
rect 8904 6780 8910 6792
rect 9125 6783 9183 6789
rect 9125 6780 9137 6783
rect 8904 6752 9137 6780
rect 8904 6740 8910 6752
rect 9125 6749 9137 6752
rect 9171 6749 9183 6783
rect 9125 6743 9183 6749
rect 9585 6783 9643 6789
rect 9585 6749 9597 6783
rect 9631 6780 9643 6783
rect 9674 6780 9680 6792
rect 9631 6752 9680 6780
rect 9631 6749 9643 6752
rect 9585 6743 9643 6749
rect 9674 6740 9680 6752
rect 9732 6740 9738 6792
rect 9766 6740 9772 6792
rect 9824 6740 9830 6792
rect 10152 6789 10180 6820
rect 12084 6820 12204 6848
rect 10137 6783 10195 6789
rect 10137 6749 10149 6783
rect 10183 6749 10195 6783
rect 10137 6743 10195 6749
rect 10318 6740 10324 6792
rect 10376 6740 10382 6792
rect 12084 6789 12112 6820
rect 12069 6783 12127 6789
rect 12069 6749 12081 6783
rect 12115 6749 12127 6783
rect 12069 6743 12127 6749
rect 12161 6783 12219 6789
rect 12161 6749 12173 6783
rect 12207 6780 12219 6783
rect 12434 6780 12440 6792
rect 12207 6752 12440 6780
rect 12207 6749 12219 6752
rect 12161 6743 12219 6749
rect 12434 6740 12440 6752
rect 12492 6740 12498 6792
rect 12544 6780 12572 6888
rect 12618 6876 12624 6928
rect 12676 6876 12682 6928
rect 14366 6876 14372 6928
rect 14424 6916 14430 6928
rect 15562 6916 15568 6928
rect 14424 6888 15568 6916
rect 14424 6876 14430 6888
rect 15562 6876 15568 6888
rect 15620 6916 15626 6928
rect 15838 6916 15844 6928
rect 15620 6888 15844 6916
rect 15620 6876 15626 6888
rect 15838 6876 15844 6888
rect 15896 6876 15902 6928
rect 12636 6848 12664 6876
rect 14182 6848 14188 6860
rect 12636 6820 12756 6848
rect 12728 6789 12756 6820
rect 13924 6820 14188 6848
rect 12621 6783 12679 6789
rect 12621 6780 12633 6783
rect 12544 6752 12633 6780
rect 12621 6749 12633 6752
rect 12667 6749 12679 6783
rect 12621 6743 12679 6749
rect 12713 6783 12771 6789
rect 12713 6749 12725 6783
rect 12759 6749 12771 6783
rect 12713 6743 12771 6749
rect 12894 6740 12900 6792
rect 12952 6740 12958 6792
rect 12986 6740 12992 6792
rect 13044 6740 13050 6792
rect 13262 6740 13268 6792
rect 13320 6740 13326 6792
rect 13541 6783 13599 6789
rect 13541 6749 13553 6783
rect 13587 6749 13599 6783
rect 13541 6743 13599 6749
rect 13633 6783 13691 6789
rect 13633 6749 13645 6783
rect 13679 6780 13691 6783
rect 13722 6780 13728 6792
rect 13679 6752 13728 6780
rect 13679 6749 13691 6752
rect 13633 6743 13691 6749
rect 8478 6712 8484 6724
rect 7668 6684 8484 6712
rect 8478 6672 8484 6684
rect 8536 6672 8542 6724
rect 11885 6715 11943 6721
rect 11885 6681 11897 6715
rect 11931 6712 11943 6715
rect 13004 6712 13032 6740
rect 13446 6712 13452 6724
rect 11931 6684 12434 6712
rect 13004 6684 13452 6712
rect 11931 6681 11943 6684
rect 11885 6675 11943 6681
rect 5994 6604 6000 6656
rect 6052 6604 6058 6656
rect 7929 6647 7987 6653
rect 7929 6613 7941 6647
rect 7975 6644 7987 6647
rect 8386 6644 8392 6656
rect 7975 6616 8392 6644
rect 7975 6613 7987 6616
rect 7929 6607 7987 6613
rect 8386 6604 8392 6616
rect 8444 6604 8450 6656
rect 8662 6604 8668 6656
rect 8720 6604 8726 6656
rect 10226 6604 10232 6656
rect 10284 6604 10290 6656
rect 12406 6644 12434 6684
rect 13446 6672 13452 6684
rect 13504 6672 13510 6724
rect 12710 6644 12716 6656
rect 12406 6616 12716 6644
rect 12710 6604 12716 6616
rect 12768 6644 12774 6656
rect 13081 6647 13139 6653
rect 13081 6644 13093 6647
rect 12768 6616 13093 6644
rect 12768 6604 12774 6616
rect 13081 6613 13093 6616
rect 13127 6613 13139 6647
rect 13556 6644 13584 6743
rect 13722 6740 13728 6752
rect 13780 6740 13786 6792
rect 13924 6789 13952 6820
rect 14182 6808 14188 6820
rect 14240 6808 14246 6860
rect 17589 6851 17647 6857
rect 14568 6820 15056 6848
rect 13909 6783 13967 6789
rect 13909 6749 13921 6783
rect 13955 6749 13967 6783
rect 13909 6743 13967 6749
rect 14274 6740 14280 6792
rect 14332 6740 14338 6792
rect 13817 6715 13875 6721
rect 13817 6681 13829 6715
rect 13863 6712 13875 6715
rect 14292 6712 14320 6740
rect 13863 6684 14320 6712
rect 13863 6681 13875 6684
rect 13817 6675 13875 6681
rect 14568 6644 14596 6820
rect 14829 6783 14887 6789
rect 14829 6780 14841 6783
rect 14660 6752 14841 6780
rect 14660 6653 14688 6752
rect 14829 6749 14841 6752
rect 14875 6749 14887 6783
rect 14829 6743 14887 6749
rect 14918 6740 14924 6792
rect 14976 6740 14982 6792
rect 15028 6712 15056 6820
rect 17589 6817 17601 6851
rect 17635 6848 17647 6851
rect 18138 6848 18144 6860
rect 17635 6820 18144 6848
rect 17635 6817 17647 6820
rect 17589 6811 17647 6817
rect 18138 6808 18144 6820
rect 18196 6808 18202 6860
rect 18966 6808 18972 6860
rect 19024 6848 19030 6860
rect 19061 6851 19119 6857
rect 19061 6848 19073 6851
rect 19024 6820 19073 6848
rect 19024 6808 19030 6820
rect 19061 6817 19073 6820
rect 19107 6817 19119 6851
rect 19061 6811 19119 6817
rect 20073 6851 20131 6857
rect 20073 6817 20085 6851
rect 20119 6848 20131 6851
rect 20346 6848 20352 6860
rect 20119 6820 20352 6848
rect 20119 6817 20131 6820
rect 20073 6811 20131 6817
rect 20346 6808 20352 6820
rect 20404 6808 20410 6860
rect 15470 6740 15476 6792
rect 15528 6740 15534 6792
rect 15733 6783 15791 6789
rect 15733 6780 15745 6783
rect 15580 6752 15745 6780
rect 15580 6712 15608 6752
rect 15733 6749 15745 6752
rect 15779 6749 15791 6783
rect 15733 6743 15791 6749
rect 15838 6740 15844 6792
rect 15896 6740 15902 6792
rect 16482 6740 16488 6792
rect 16540 6780 16546 6792
rect 17313 6783 17371 6789
rect 17313 6780 17325 6783
rect 16540 6752 17325 6780
rect 16540 6740 16546 6752
rect 17313 6749 17325 6752
rect 17359 6749 17371 6783
rect 17313 6743 17371 6749
rect 18690 6740 18696 6792
rect 18748 6740 18754 6792
rect 21450 6740 21456 6792
rect 21508 6740 21514 6792
rect 23382 6740 23388 6792
rect 23440 6780 23446 6792
rect 23661 6783 23719 6789
rect 23661 6780 23673 6783
rect 23440 6752 23673 6780
rect 23440 6740 23446 6752
rect 23661 6749 23673 6752
rect 23707 6749 23719 6783
rect 23661 6743 23719 6749
rect 24029 6783 24087 6789
rect 24029 6749 24041 6783
rect 24075 6780 24087 6783
rect 24302 6780 24308 6792
rect 24075 6752 24308 6780
rect 24075 6749 24087 6752
rect 24029 6743 24087 6749
rect 24302 6740 24308 6752
rect 24360 6740 24366 6792
rect 15028 6684 15608 6712
rect 13556 6616 14596 6644
rect 14645 6647 14703 6653
rect 13081 6607 13139 6613
rect 14645 6613 14657 6647
rect 14691 6613 14703 6647
rect 15580 6644 15608 6684
rect 15657 6715 15715 6721
rect 15657 6681 15669 6715
rect 15703 6712 15715 6715
rect 16206 6712 16212 6724
rect 15703 6684 16212 6712
rect 15703 6681 15715 6684
rect 15657 6675 15715 6681
rect 16206 6672 16212 6684
rect 16264 6672 16270 6724
rect 16298 6644 16304 6656
rect 15580 6616 16304 6644
rect 14645 6607 14703 6613
rect 16298 6604 16304 6616
rect 16356 6604 16362 6656
rect 1104 6554 28152 6576
rect 1104 6502 4874 6554
rect 4926 6502 4938 6554
rect 4990 6502 5002 6554
rect 5054 6502 5066 6554
rect 5118 6502 5130 6554
rect 5182 6502 28152 6554
rect 1104 6480 28152 6502
rect 12526 6440 12532 6452
rect 11532 6412 12532 6440
rect 5994 6264 6000 6316
rect 6052 6304 6058 6316
rect 8021 6307 8079 6313
rect 8021 6304 8033 6307
rect 6052 6276 8033 6304
rect 6052 6264 6058 6276
rect 8021 6273 8033 6276
rect 8067 6304 8079 6307
rect 8570 6304 8576 6316
rect 8067 6276 8576 6304
rect 8067 6273 8079 6276
rect 8021 6267 8079 6273
rect 8570 6264 8576 6276
rect 8628 6264 8634 6316
rect 8938 6264 8944 6316
rect 8996 6304 9002 6316
rect 10226 6304 10232 6316
rect 8996 6276 10232 6304
rect 8996 6264 9002 6276
rect 10226 6264 10232 6276
rect 10284 6264 10290 6316
rect 11532 6313 11560 6412
rect 12526 6400 12532 6412
rect 12584 6440 12590 6452
rect 12584 6412 16344 6440
rect 12584 6400 12590 6412
rect 11793 6375 11851 6381
rect 11793 6341 11805 6375
rect 11839 6372 11851 6375
rect 11882 6372 11888 6384
rect 11839 6344 11888 6372
rect 11839 6341 11851 6344
rect 11793 6335 11851 6341
rect 11882 6332 11888 6344
rect 11940 6332 11946 6384
rect 13170 6372 13176 6384
rect 13018 6344 13176 6372
rect 13170 6332 13176 6344
rect 13228 6372 13234 6384
rect 13228 6344 14780 6372
rect 13228 6332 13234 6344
rect 11517 6307 11575 6313
rect 11517 6273 11529 6307
rect 11563 6273 11575 6307
rect 11517 6267 11575 6273
rect 13446 6264 13452 6316
rect 13504 6264 13510 6316
rect 13541 6307 13599 6313
rect 13541 6273 13553 6307
rect 13587 6304 13599 6307
rect 13722 6304 13728 6316
rect 13587 6276 13728 6304
rect 13587 6273 13599 6276
rect 13541 6267 13599 6273
rect 8113 6239 8171 6245
rect 8113 6205 8125 6239
rect 8159 6205 8171 6239
rect 8113 6199 8171 6205
rect 8128 6168 8156 6199
rect 8386 6196 8392 6248
rect 8444 6236 8450 6248
rect 8849 6239 8907 6245
rect 8849 6236 8861 6239
rect 8444 6208 8861 6236
rect 8444 6196 8450 6208
rect 8849 6205 8861 6208
rect 8895 6205 8907 6239
rect 8849 6199 8907 6205
rect 9309 6239 9367 6245
rect 9309 6205 9321 6239
rect 9355 6236 9367 6239
rect 9674 6236 9680 6248
rect 9355 6208 9680 6236
rect 9355 6205 9367 6208
rect 9309 6199 9367 6205
rect 9674 6196 9680 6208
rect 9732 6196 9738 6248
rect 10318 6196 10324 6248
rect 10376 6236 10382 6248
rect 13265 6239 13323 6245
rect 10376 6208 13216 6236
rect 10376 6196 10382 6208
rect 8754 6168 8760 6180
rect 8128 6140 8760 6168
rect 8754 6128 8760 6140
rect 8812 6128 8818 6180
rect 13188 6168 13216 6208
rect 13265 6205 13277 6239
rect 13311 6236 13323 6239
rect 13556 6236 13584 6267
rect 13722 6264 13728 6276
rect 13780 6264 13786 6316
rect 13311 6208 13584 6236
rect 13311 6205 13323 6208
rect 13265 6199 13323 6205
rect 14274 6196 14280 6248
rect 14332 6236 14338 6248
rect 14553 6239 14611 6245
rect 14553 6236 14565 6239
rect 14332 6208 14565 6236
rect 14332 6196 14338 6208
rect 14553 6205 14565 6208
rect 14599 6205 14611 6239
rect 14752 6236 14780 6344
rect 16022 6332 16028 6384
rect 16080 6332 16086 6384
rect 16316 6313 16344 6412
rect 18598 6400 18604 6452
rect 18656 6400 18662 6452
rect 27614 6400 27620 6452
rect 27672 6400 27678 6452
rect 17034 6332 17040 6384
rect 17092 6372 17098 6384
rect 17129 6375 17187 6381
rect 17129 6372 17141 6375
rect 17092 6344 17141 6372
rect 17092 6332 17098 6344
rect 17129 6341 17141 6344
rect 17175 6341 17187 6375
rect 18690 6372 18696 6384
rect 18354 6358 18696 6372
rect 17129 6335 17187 6341
rect 18340 6344 18696 6358
rect 16301 6307 16359 6313
rect 14936 6236 14964 6290
rect 16301 6273 16313 6307
rect 16347 6304 16359 6307
rect 16482 6304 16488 6316
rect 16347 6276 16488 6304
rect 16347 6273 16359 6276
rect 16301 6267 16359 6273
rect 16482 6264 16488 6276
rect 16540 6304 16546 6316
rect 16853 6307 16911 6313
rect 16853 6304 16865 6307
rect 16540 6276 16865 6304
rect 16540 6264 16546 6276
rect 16853 6273 16865 6276
rect 16899 6273 16911 6307
rect 16853 6267 16911 6273
rect 18340 6236 18368 6344
rect 18690 6332 18696 6344
rect 18748 6332 18754 6384
rect 27798 6264 27804 6316
rect 27856 6264 27862 6316
rect 14752 6208 18368 6236
rect 14553 6199 14611 6205
rect 13814 6168 13820 6180
rect 13188 6140 13820 6168
rect 13814 6128 13820 6140
rect 13872 6128 13878 6180
rect 1104 6010 28152 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 28152 6010
rect 1104 5936 28152 5958
rect 8478 5856 8484 5908
rect 8536 5896 8542 5908
rect 8665 5899 8723 5905
rect 8665 5896 8677 5899
rect 8536 5868 8677 5896
rect 8536 5856 8542 5868
rect 8665 5865 8677 5868
rect 8711 5865 8723 5899
rect 8665 5859 8723 5865
rect 13262 5856 13268 5908
rect 13320 5896 13326 5908
rect 15470 5896 15476 5908
rect 13320 5868 15476 5896
rect 13320 5856 13326 5868
rect 15470 5856 15476 5868
rect 15528 5856 15534 5908
rect 27617 5899 27675 5905
rect 27617 5865 27629 5899
rect 27663 5896 27675 5899
rect 27706 5896 27712 5908
rect 27663 5868 27712 5896
rect 27663 5865 27675 5868
rect 27617 5859 27675 5865
rect 27706 5856 27712 5868
rect 27764 5856 27770 5908
rect 8938 5760 8944 5772
rect 8496 5732 8944 5760
rect 8386 5652 8392 5704
rect 8444 5652 8450 5704
rect 8496 5701 8524 5732
rect 8938 5720 8944 5732
rect 8996 5720 9002 5772
rect 8481 5695 8539 5701
rect 8481 5661 8493 5695
rect 8527 5661 8539 5695
rect 8481 5655 8539 5661
rect 8662 5652 8668 5704
rect 8720 5652 8726 5704
rect 27798 5652 27804 5704
rect 27856 5652 27862 5704
rect 1104 5466 28152 5488
rect 1104 5414 4874 5466
rect 4926 5414 4938 5466
rect 4990 5414 5002 5466
rect 5054 5414 5066 5466
rect 5118 5414 5130 5466
rect 5182 5414 28152 5466
rect 1104 5392 28152 5414
rect 1104 4922 28152 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 28152 4922
rect 1104 4848 28152 4870
rect 1104 4378 28152 4400
rect 1104 4326 4874 4378
rect 4926 4326 4938 4378
rect 4990 4326 5002 4378
rect 5054 4326 5066 4378
rect 5118 4326 5130 4378
rect 5182 4326 28152 4378
rect 1104 4304 28152 4326
rect 1104 3834 28152 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 28152 3834
rect 1104 3760 28152 3782
rect 1104 3290 28152 3312
rect 1104 3238 4874 3290
rect 4926 3238 4938 3290
rect 4990 3238 5002 3290
rect 5054 3238 5066 3290
rect 5118 3238 5130 3290
rect 5182 3238 28152 3290
rect 1104 3216 28152 3238
rect 1104 2746 28152 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 28152 2746
rect 1104 2672 28152 2694
rect 6086 2592 6092 2644
rect 6144 2592 6150 2644
rect 9306 2592 9312 2644
rect 9364 2592 9370 2644
rect 5810 2388 5816 2440
rect 5868 2428 5874 2440
rect 5905 2431 5963 2437
rect 5905 2428 5917 2431
rect 5868 2400 5917 2428
rect 5868 2388 5874 2400
rect 5905 2397 5917 2400
rect 5951 2397 5963 2431
rect 5905 2391 5963 2397
rect 9030 2388 9036 2440
rect 9088 2428 9094 2440
rect 9125 2431 9183 2437
rect 9125 2428 9137 2431
rect 9088 2400 9137 2428
rect 9088 2388 9094 2400
rect 9125 2397 9137 2400
rect 9171 2397 9183 2431
rect 9125 2391 9183 2397
rect 1104 2202 28152 2224
rect 1104 2150 4874 2202
rect 4926 2150 4938 2202
rect 4990 2150 5002 2202
rect 5054 2150 5066 2202
rect 5118 2150 5130 2202
rect 5182 2150 28152 2202
rect 1104 2128 28152 2150
<< via1 >>
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 11796 28747 11848 28756
rect 11796 28713 11805 28747
rect 11805 28713 11839 28747
rect 11839 28713 11848 28747
rect 11796 28704 11848 28713
rect 12348 28704 12400 28756
rect 13084 28747 13136 28756
rect 13084 28713 13093 28747
rect 13093 28713 13127 28747
rect 13127 28713 13136 28747
rect 13084 28704 13136 28713
rect 13728 28747 13780 28756
rect 13728 28713 13737 28747
rect 13737 28713 13771 28747
rect 13771 28713 13780 28747
rect 13728 28704 13780 28713
rect 14372 28747 14424 28756
rect 14372 28713 14381 28747
rect 14381 28713 14415 28747
rect 14415 28713 14424 28747
rect 14372 28704 14424 28713
rect 15016 28747 15068 28756
rect 15016 28713 15025 28747
rect 15025 28713 15059 28747
rect 15059 28713 15068 28747
rect 15016 28704 15068 28713
rect 15660 28747 15712 28756
rect 15660 28713 15669 28747
rect 15669 28713 15703 28747
rect 15703 28713 15712 28747
rect 15660 28704 15712 28713
rect 16304 28747 16356 28756
rect 16304 28713 16313 28747
rect 16313 28713 16347 28747
rect 16347 28713 16356 28747
rect 16304 28704 16356 28713
rect 16948 28747 17000 28756
rect 16948 28713 16957 28747
rect 16957 28713 16991 28747
rect 16991 28713 17000 28747
rect 16948 28704 17000 28713
rect 17592 28747 17644 28756
rect 17592 28713 17601 28747
rect 17601 28713 17635 28747
rect 17635 28713 17644 28747
rect 17592 28704 17644 28713
rect 18236 28747 18288 28756
rect 18236 28713 18245 28747
rect 18245 28713 18279 28747
rect 18279 28713 18288 28747
rect 18236 28704 18288 28713
rect 18880 28747 18932 28756
rect 18880 28713 18889 28747
rect 18889 28713 18923 28747
rect 18923 28713 18932 28747
rect 18880 28704 18932 28713
rect 19616 28747 19668 28756
rect 19616 28713 19625 28747
rect 19625 28713 19659 28747
rect 19659 28713 19668 28747
rect 19616 28704 19668 28713
rect 20260 28747 20312 28756
rect 20260 28713 20269 28747
rect 20269 28713 20303 28747
rect 20303 28713 20312 28747
rect 20260 28704 20312 28713
rect 20536 28704 20588 28756
rect 21548 28747 21600 28756
rect 21548 28713 21557 28747
rect 21557 28713 21591 28747
rect 21591 28713 21600 28747
rect 21548 28704 21600 28713
rect 22008 28704 22060 28756
rect 22836 28747 22888 28756
rect 22836 28713 22845 28747
rect 22845 28713 22879 28747
rect 22879 28713 22888 28747
rect 22836 28704 22888 28713
rect 23388 28704 23440 28756
rect 24124 28747 24176 28756
rect 24124 28713 24133 28747
rect 24133 28713 24167 28747
rect 24167 28713 24176 28747
rect 24124 28704 24176 28713
rect 24768 28747 24820 28756
rect 24768 28713 24777 28747
rect 24777 28713 24811 28747
rect 24811 28713 24820 28747
rect 24768 28704 24820 28713
rect 25412 28747 25464 28756
rect 25412 28713 25421 28747
rect 25421 28713 25455 28747
rect 25455 28713 25464 28747
rect 25412 28704 25464 28713
rect 26056 28747 26108 28756
rect 26056 28713 26065 28747
rect 26065 28713 26099 28747
rect 26099 28713 26108 28747
rect 26056 28704 26108 28713
rect 26700 28747 26752 28756
rect 26700 28713 26709 28747
rect 26709 28713 26743 28747
rect 26743 28713 26752 28747
rect 26700 28704 26752 28713
rect 27344 28747 27396 28756
rect 27344 28713 27353 28747
rect 27353 28713 27387 28747
rect 27387 28713 27396 28747
rect 27344 28704 27396 28713
rect 27804 28704 27856 28756
rect 11980 28543 12032 28552
rect 11980 28509 11989 28543
rect 11989 28509 12023 28543
rect 12023 28509 12032 28543
rect 11980 28500 12032 28509
rect 13268 28543 13320 28552
rect 13268 28509 13277 28543
rect 13277 28509 13311 28543
rect 13311 28509 13320 28543
rect 13268 28500 13320 28509
rect 18144 28636 18196 28688
rect 17960 28568 18012 28620
rect 15844 28543 15896 28552
rect 15844 28509 15853 28543
rect 15853 28509 15887 28543
rect 15887 28509 15896 28543
rect 15844 28500 15896 28509
rect 16948 28500 17000 28552
rect 17132 28543 17184 28552
rect 17132 28509 17141 28543
rect 17141 28509 17175 28543
rect 17175 28509 17184 28543
rect 17132 28500 17184 28509
rect 17868 28500 17920 28552
rect 17408 28432 17460 28484
rect 19984 28568 20036 28620
rect 19064 28543 19116 28552
rect 19064 28509 19073 28543
rect 19073 28509 19107 28543
rect 19107 28509 19116 28543
rect 19064 28500 19116 28509
rect 19432 28543 19484 28552
rect 19432 28509 19441 28543
rect 19441 28509 19475 28543
rect 19475 28509 19484 28543
rect 19432 28500 19484 28509
rect 19892 28500 19944 28552
rect 20444 28500 20496 28552
rect 21364 28543 21416 28552
rect 21364 28509 21373 28543
rect 21373 28509 21407 28543
rect 21407 28509 21416 28543
rect 21364 28500 21416 28509
rect 22284 28543 22336 28552
rect 22284 28509 22293 28543
rect 22293 28509 22327 28543
rect 22327 28509 22336 28543
rect 22284 28500 22336 28509
rect 22652 28543 22704 28552
rect 22652 28509 22661 28543
rect 22661 28509 22695 28543
rect 22695 28509 22704 28543
rect 22652 28500 22704 28509
rect 23296 28543 23348 28552
rect 23296 28509 23305 28543
rect 23305 28509 23339 28543
rect 23339 28509 23348 28543
rect 23296 28500 23348 28509
rect 23940 28543 23992 28552
rect 23940 28509 23949 28543
rect 23949 28509 23983 28543
rect 23983 28509 23992 28543
rect 23940 28500 23992 28509
rect 24584 28543 24636 28552
rect 24584 28509 24593 28543
rect 24593 28509 24627 28543
rect 24627 28509 24636 28543
rect 24584 28500 24636 28509
rect 24952 28500 25004 28552
rect 25872 28543 25924 28552
rect 25872 28509 25881 28543
rect 25881 28509 25915 28543
rect 25915 28509 25924 28543
rect 25872 28500 25924 28509
rect 26056 28500 26108 28552
rect 26792 28500 26844 28552
rect 21456 28432 21508 28484
rect 26148 28432 26200 28484
rect 17224 28364 17276 28416
rect 17776 28364 17828 28416
rect 18696 28364 18748 28416
rect 20076 28364 20128 28416
rect 4874 28262 4926 28314
rect 4938 28262 4990 28314
rect 5002 28262 5054 28314
rect 5066 28262 5118 28314
rect 5130 28262 5182 28314
rect 17132 28160 17184 28212
rect 19064 28160 19116 28212
rect 20444 28203 20496 28212
rect 20444 28169 20453 28203
rect 20453 28169 20487 28203
rect 20487 28169 20496 28203
rect 20444 28160 20496 28169
rect 24952 28203 25004 28212
rect 24952 28169 24961 28203
rect 24961 28169 24995 28203
rect 24995 28169 25004 28203
rect 24952 28160 25004 28169
rect 28724 28160 28776 28212
rect 7472 27956 7524 28008
rect 11060 28067 11112 28076
rect 13268 28092 13320 28144
rect 11060 28033 11099 28067
rect 11099 28033 11112 28067
rect 11060 28024 11112 28033
rect 11704 28024 11756 28076
rect 11980 28024 12032 28076
rect 18604 28024 18656 28076
rect 18696 28067 18748 28076
rect 18696 28033 18705 28067
rect 18705 28033 18739 28067
rect 18739 28033 18748 28067
rect 18696 28024 18748 28033
rect 15844 27956 15896 28008
rect 19064 27956 19116 28008
rect 19524 28024 19576 28076
rect 19616 27956 19668 28008
rect 10692 27931 10744 27940
rect 10692 27897 10701 27931
rect 10701 27897 10735 27931
rect 10735 27897 10744 27931
rect 10692 27888 10744 27897
rect 11152 27888 11204 27940
rect 18052 27888 18104 27940
rect 19156 27888 19208 27940
rect 19708 27888 19760 27940
rect 20076 28067 20128 28076
rect 20076 28033 20091 28067
rect 20091 28033 20125 28067
rect 20125 28033 20128 28067
rect 20076 28024 20128 28033
rect 19984 27999 20036 28008
rect 19984 27965 19993 27999
rect 19993 27965 20027 27999
rect 20027 27965 20036 27999
rect 19984 27956 20036 27965
rect 20352 28067 20404 28076
rect 20352 28033 20361 28067
rect 20361 28033 20395 28067
rect 20395 28033 20404 28067
rect 20352 28024 20404 28033
rect 21088 27956 21140 28008
rect 20996 27888 21048 27940
rect 21640 28067 21692 28076
rect 21640 28033 21649 28067
rect 21649 28033 21683 28067
rect 21683 28033 21692 28067
rect 21640 28024 21692 28033
rect 22100 28024 22152 28076
rect 23388 28024 23440 28076
rect 24952 28024 25004 28076
rect 25044 28067 25096 28076
rect 25044 28033 25053 28067
rect 25053 28033 25087 28067
rect 25087 28033 25096 28067
rect 25044 28024 25096 28033
rect 27160 28067 27212 28076
rect 27160 28033 27169 28067
rect 27169 28033 27203 28067
rect 27203 28033 27212 28067
rect 27160 28024 27212 28033
rect 22376 27956 22428 28008
rect 25412 27956 25464 28008
rect 24032 27888 24084 27940
rect 26240 27888 26292 27940
rect 27988 27888 28040 27940
rect 11244 27820 11296 27872
rect 18788 27820 18840 27872
rect 21548 27863 21600 27872
rect 21548 27829 21557 27863
rect 21557 27829 21591 27863
rect 21591 27829 21600 27863
rect 21548 27820 21600 27829
rect 22100 27820 22152 27872
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 2780 27616 2832 27668
rect 3148 27548 3200 27600
rect 4620 27480 4672 27532
rect 5448 27548 5500 27600
rect 5724 27480 5776 27532
rect 2044 27412 2096 27464
rect 5172 27412 5224 27464
rect 5908 27412 5960 27464
rect 6000 27455 6052 27464
rect 6000 27421 6009 27455
rect 6009 27421 6043 27455
rect 6043 27421 6052 27455
rect 6000 27412 6052 27421
rect 5632 27344 5684 27396
rect 5724 27344 5776 27396
rect 6184 27455 6236 27464
rect 6184 27421 6193 27455
rect 6193 27421 6227 27455
rect 6227 27421 6236 27455
rect 6184 27412 6236 27421
rect 6920 27616 6972 27668
rect 10324 27659 10376 27668
rect 10324 27625 10333 27659
rect 10333 27625 10367 27659
rect 10367 27625 10376 27659
rect 10324 27616 10376 27625
rect 6736 27548 6788 27600
rect 7472 27548 7524 27600
rect 10508 27548 10560 27600
rect 11060 27616 11112 27668
rect 10968 27548 11020 27600
rect 6828 27412 6880 27464
rect 7472 27455 7524 27464
rect 7472 27421 7481 27455
rect 7481 27421 7515 27455
rect 7515 27421 7524 27455
rect 7472 27412 7524 27421
rect 7656 27455 7708 27464
rect 7656 27421 7665 27455
rect 7665 27421 7699 27455
rect 7699 27421 7708 27455
rect 7656 27412 7708 27421
rect 10600 27455 10652 27464
rect 10600 27421 10609 27455
rect 10609 27421 10643 27455
rect 10643 27421 10652 27455
rect 10600 27412 10652 27421
rect 10784 27455 10836 27464
rect 10784 27421 10793 27455
rect 10793 27421 10827 27455
rect 10827 27421 10836 27455
rect 10784 27412 10836 27421
rect 11244 27412 11296 27464
rect 16948 27591 17000 27600
rect 16948 27557 16957 27591
rect 16957 27557 16991 27591
rect 16991 27557 17000 27591
rect 16948 27548 17000 27557
rect 17224 27591 17276 27600
rect 17224 27557 17233 27591
rect 17233 27557 17267 27591
rect 17267 27557 17276 27591
rect 17224 27548 17276 27557
rect 17776 27548 17828 27600
rect 18236 27616 18288 27668
rect 18788 27659 18840 27668
rect 18788 27625 18797 27659
rect 18797 27625 18831 27659
rect 18831 27625 18840 27659
rect 18788 27616 18840 27625
rect 19248 27616 19300 27668
rect 19892 27659 19944 27668
rect 19892 27625 19901 27659
rect 19901 27625 19935 27659
rect 19935 27625 19944 27659
rect 19892 27616 19944 27625
rect 20076 27659 20128 27668
rect 20076 27625 20085 27659
rect 20085 27625 20119 27659
rect 20119 27625 20128 27659
rect 20076 27616 20128 27625
rect 20812 27659 20864 27668
rect 20812 27625 20821 27659
rect 20821 27625 20855 27659
rect 20855 27625 20864 27659
rect 20812 27616 20864 27625
rect 18604 27591 18656 27600
rect 18604 27557 18613 27591
rect 18613 27557 18647 27591
rect 18647 27557 18656 27591
rect 18604 27548 18656 27557
rect 21088 27591 21140 27600
rect 21088 27557 21097 27591
rect 21097 27557 21131 27591
rect 21131 27557 21140 27591
rect 21088 27548 21140 27557
rect 11704 27455 11756 27464
rect 11704 27421 11743 27455
rect 11743 27421 11756 27455
rect 11704 27412 11756 27421
rect 11888 27455 11940 27464
rect 11888 27421 11897 27455
rect 11897 27421 11931 27455
rect 11931 27421 11940 27455
rect 11888 27412 11940 27421
rect 16948 27455 17000 27464
rect 16948 27421 16957 27455
rect 16957 27421 16991 27455
rect 16991 27421 17000 27455
rect 16948 27412 17000 27421
rect 18696 27480 18748 27532
rect 18788 27480 18840 27532
rect 18512 27455 18564 27464
rect 5356 27276 5408 27328
rect 5448 27319 5500 27328
rect 5448 27285 5457 27319
rect 5457 27285 5491 27319
rect 5491 27285 5500 27319
rect 5448 27276 5500 27285
rect 5540 27276 5592 27328
rect 18512 27421 18521 27455
rect 18521 27421 18555 27455
rect 18555 27421 18564 27455
rect 18512 27412 18564 27421
rect 19248 27412 19300 27464
rect 19616 27412 19668 27464
rect 20260 27412 20312 27464
rect 6736 27276 6788 27328
rect 6828 27276 6880 27328
rect 19156 27344 19208 27396
rect 10324 27276 10376 27328
rect 10416 27276 10468 27328
rect 10600 27276 10652 27328
rect 11980 27276 12032 27328
rect 17960 27319 18012 27328
rect 17960 27285 17969 27319
rect 17969 27285 18003 27319
rect 18003 27285 18012 27319
rect 17960 27276 18012 27285
rect 18236 27276 18288 27328
rect 18328 27276 18380 27328
rect 19064 27276 19116 27328
rect 19524 27276 19576 27328
rect 19800 27387 19852 27396
rect 19800 27353 19809 27387
rect 19809 27353 19843 27387
rect 19843 27353 19852 27387
rect 19800 27344 19852 27353
rect 20168 27344 20220 27396
rect 20904 27455 20956 27464
rect 20904 27421 20913 27455
rect 20913 27421 20947 27455
rect 20947 27421 20956 27455
rect 20904 27412 20956 27421
rect 21364 27659 21416 27668
rect 21364 27625 21373 27659
rect 21373 27625 21407 27659
rect 21407 27625 21416 27659
rect 21364 27616 21416 27625
rect 22284 27616 22336 27668
rect 23940 27616 23992 27668
rect 24584 27616 24636 27668
rect 24676 27616 24728 27668
rect 25044 27616 25096 27668
rect 21456 27591 21508 27600
rect 21456 27557 21465 27591
rect 21465 27557 21499 27591
rect 21499 27557 21508 27591
rect 21456 27548 21508 27557
rect 22560 27548 22612 27600
rect 25964 27616 26016 27668
rect 26792 27659 26844 27668
rect 26792 27625 26801 27659
rect 26801 27625 26835 27659
rect 26835 27625 26844 27659
rect 26792 27616 26844 27625
rect 27160 27616 27212 27668
rect 21640 27480 21692 27532
rect 22100 27480 22152 27532
rect 24860 27480 24912 27532
rect 25320 27523 25372 27532
rect 25320 27489 25345 27523
rect 25345 27489 25372 27523
rect 25320 27480 25372 27489
rect 25780 27548 25832 27600
rect 20996 27344 21048 27396
rect 22192 27387 22244 27396
rect 22192 27353 22201 27387
rect 22201 27353 22235 27387
rect 22235 27353 22244 27387
rect 22192 27344 22244 27353
rect 22560 27387 22612 27396
rect 22560 27353 22578 27387
rect 22578 27353 22612 27387
rect 22560 27344 22612 27353
rect 23020 27455 23072 27464
rect 23020 27421 23029 27455
rect 23029 27421 23063 27455
rect 23063 27421 23072 27455
rect 23020 27412 23072 27421
rect 23112 27455 23164 27464
rect 23112 27421 23121 27455
rect 23121 27421 23155 27455
rect 23155 27421 23164 27455
rect 23112 27412 23164 27421
rect 23388 27455 23440 27464
rect 23388 27421 23397 27455
rect 23397 27421 23431 27455
rect 23431 27421 23440 27455
rect 23388 27412 23440 27421
rect 24032 27455 24084 27464
rect 24032 27421 24041 27455
rect 24041 27421 24075 27455
rect 24075 27421 24084 27455
rect 24032 27412 24084 27421
rect 24216 27455 24268 27464
rect 24216 27421 24225 27455
rect 24225 27421 24259 27455
rect 24259 27421 24268 27455
rect 24216 27412 24268 27421
rect 24400 27412 24452 27464
rect 20812 27276 20864 27328
rect 22928 27276 22980 27328
rect 23756 27344 23808 27396
rect 24676 27412 24728 27464
rect 25504 27412 25556 27464
rect 25780 27455 25832 27464
rect 25780 27421 25789 27455
rect 25789 27421 25823 27455
rect 25823 27421 25832 27455
rect 25780 27412 25832 27421
rect 25964 27412 26016 27464
rect 26332 27523 26384 27532
rect 26332 27489 26341 27523
rect 26341 27489 26375 27523
rect 26375 27489 26384 27523
rect 26332 27480 26384 27489
rect 26240 27344 26292 27396
rect 26792 27455 26844 27464
rect 26792 27421 26801 27455
rect 26801 27421 26835 27455
rect 26835 27421 26844 27455
rect 26792 27412 26844 27421
rect 25780 27276 25832 27328
rect 25964 27319 26016 27328
rect 25964 27285 25973 27319
rect 25973 27285 26007 27319
rect 26007 27285 26016 27319
rect 25964 27276 26016 27285
rect 4874 27174 4926 27226
rect 4938 27174 4990 27226
rect 5002 27174 5054 27226
rect 5066 27174 5118 27226
rect 5130 27174 5182 27226
rect 5264 27072 5316 27124
rect 2780 27047 2832 27056
rect 2780 27013 2789 27047
rect 2789 27013 2823 27047
rect 2823 27013 2832 27047
rect 2780 27004 2832 27013
rect 2044 26936 2096 26988
rect 3516 26979 3568 26988
rect 3516 26945 3525 26979
rect 3525 26945 3559 26979
rect 3559 26945 3568 26979
rect 3516 26936 3568 26945
rect 5448 27004 5500 27056
rect 6644 27004 6696 27056
rect 2136 26911 2188 26920
rect 2136 26877 2145 26911
rect 2145 26877 2179 26911
rect 2179 26877 2188 26911
rect 2136 26868 2188 26877
rect 2596 26911 2648 26920
rect 2596 26877 2605 26911
rect 2605 26877 2639 26911
rect 2639 26877 2648 26911
rect 2596 26868 2648 26877
rect 3056 26800 3108 26852
rect 2504 26732 2556 26784
rect 3792 26868 3844 26920
rect 3884 26911 3936 26920
rect 3884 26877 3893 26911
rect 3893 26877 3927 26911
rect 3927 26877 3936 26911
rect 3884 26868 3936 26877
rect 5540 26979 5592 26988
rect 5540 26945 5549 26979
rect 5549 26945 5583 26979
rect 5583 26945 5592 26979
rect 5540 26936 5592 26945
rect 6552 26979 6604 26988
rect 6552 26945 6561 26979
rect 6561 26945 6595 26979
rect 6595 26945 6604 26979
rect 6552 26936 6604 26945
rect 6920 26936 6972 26988
rect 7656 27004 7708 27056
rect 11060 27072 11112 27124
rect 11980 27047 12032 27056
rect 11980 27013 11989 27047
rect 11989 27013 12023 27047
rect 12023 27013 12032 27047
rect 11980 27004 12032 27013
rect 12348 27072 12400 27124
rect 17408 27115 17460 27124
rect 17408 27081 17417 27115
rect 17417 27081 17451 27115
rect 17451 27081 17460 27115
rect 17408 27072 17460 27081
rect 18052 27072 18104 27124
rect 18144 27115 18196 27124
rect 18144 27081 18153 27115
rect 18153 27081 18187 27115
rect 18187 27081 18196 27115
rect 18144 27072 18196 27081
rect 9128 26979 9180 26988
rect 9128 26945 9137 26979
rect 9137 26945 9171 26979
rect 9171 26945 9180 26979
rect 9128 26936 9180 26945
rect 10600 26936 10652 26988
rect 10784 26979 10836 26988
rect 10784 26945 10793 26979
rect 10793 26945 10827 26979
rect 10827 26945 10836 26979
rect 10784 26936 10836 26945
rect 10968 26979 11020 26988
rect 10968 26945 10977 26979
rect 10977 26945 11011 26979
rect 11011 26945 11020 26979
rect 10968 26936 11020 26945
rect 11060 26936 11112 26988
rect 12992 27004 13044 27056
rect 16948 27004 17000 27056
rect 12716 26979 12768 26988
rect 12716 26945 12725 26979
rect 12725 26945 12759 26979
rect 12759 26945 12768 26979
rect 12716 26936 12768 26945
rect 4804 26911 4856 26920
rect 4804 26877 4813 26911
rect 4813 26877 4847 26911
rect 4847 26877 4856 26911
rect 4804 26868 4856 26877
rect 5448 26911 5500 26920
rect 5448 26877 5457 26911
rect 5457 26877 5491 26911
rect 5491 26877 5500 26911
rect 5448 26868 5500 26877
rect 5724 26911 5776 26920
rect 5724 26877 5733 26911
rect 5733 26877 5767 26911
rect 5767 26877 5776 26911
rect 5724 26868 5776 26877
rect 6828 26868 6880 26920
rect 5816 26843 5868 26852
rect 5816 26809 5825 26843
rect 5825 26809 5859 26843
rect 5859 26809 5868 26843
rect 5816 26800 5868 26809
rect 5908 26800 5960 26852
rect 7012 26800 7064 26852
rect 9864 26911 9916 26920
rect 9864 26877 9873 26911
rect 9873 26877 9907 26911
rect 9907 26877 9916 26911
rect 9864 26868 9916 26877
rect 17960 26936 18012 26988
rect 18512 27047 18564 27056
rect 18512 27013 18521 27047
rect 18521 27013 18555 27047
rect 18555 27013 18564 27047
rect 18512 27004 18564 27013
rect 19432 27072 19484 27124
rect 20352 27072 20404 27124
rect 20996 27115 21048 27124
rect 20996 27081 21005 27115
rect 21005 27081 21039 27115
rect 21039 27081 21048 27115
rect 20996 27072 21048 27081
rect 21548 27072 21600 27124
rect 22652 27072 22704 27124
rect 23296 27072 23348 27124
rect 24216 27072 24268 27124
rect 24768 27115 24820 27124
rect 24768 27081 24777 27115
rect 24777 27081 24811 27115
rect 24811 27081 24820 27115
rect 24768 27072 24820 27081
rect 25872 27072 25924 27124
rect 26056 27072 26108 27124
rect 18696 26936 18748 26988
rect 4712 26732 4764 26784
rect 4988 26732 5040 26784
rect 5632 26732 5684 26784
rect 6184 26732 6236 26784
rect 6828 26775 6880 26784
rect 6828 26741 6837 26775
rect 6837 26741 6871 26775
rect 6871 26741 6880 26775
rect 6828 26732 6880 26741
rect 6920 26775 6972 26784
rect 6920 26741 6929 26775
rect 6929 26741 6963 26775
rect 6963 26741 6972 26775
rect 6920 26732 6972 26741
rect 9956 26800 10008 26852
rect 10416 26800 10468 26852
rect 7656 26732 7708 26784
rect 8760 26732 8812 26784
rect 9772 26732 9824 26784
rect 10232 26732 10284 26784
rect 10600 26732 10652 26784
rect 17868 26843 17920 26852
rect 17868 26809 17877 26843
rect 17877 26809 17911 26843
rect 17911 26809 17920 26843
rect 17868 26800 17920 26809
rect 17960 26800 18012 26852
rect 18788 26800 18840 26852
rect 19524 26979 19576 26988
rect 19524 26945 19533 26979
rect 19533 26945 19567 26979
rect 19567 26945 19576 26979
rect 19984 27004 20036 27056
rect 19524 26936 19576 26945
rect 19800 26979 19852 26988
rect 19800 26945 19809 26979
rect 19809 26945 19843 26979
rect 19843 26945 19852 26979
rect 19800 26936 19852 26945
rect 11244 26732 11296 26784
rect 11520 26775 11572 26784
rect 11520 26741 11529 26775
rect 11529 26741 11563 26775
rect 11563 26741 11572 26775
rect 11520 26732 11572 26741
rect 11704 26775 11756 26784
rect 11704 26741 11713 26775
rect 11713 26741 11747 26775
rect 11747 26741 11756 26775
rect 11704 26732 11756 26741
rect 12532 26732 12584 26784
rect 18328 26775 18380 26784
rect 18328 26741 18337 26775
rect 18337 26741 18371 26775
rect 18371 26741 18380 26775
rect 18328 26732 18380 26741
rect 18512 26732 18564 26784
rect 19984 26911 20036 26920
rect 19984 26877 19993 26911
rect 19993 26877 20027 26911
rect 20027 26877 20036 26911
rect 19984 26868 20036 26877
rect 20260 26979 20312 26988
rect 20260 26945 20269 26979
rect 20269 26945 20303 26979
rect 20303 26945 20312 26979
rect 20260 26936 20312 26945
rect 20904 27004 20956 27056
rect 20444 26868 20496 26920
rect 19248 26800 19300 26852
rect 20628 26936 20680 26988
rect 20996 26936 21048 26988
rect 21916 27004 21968 27056
rect 22284 27004 22336 27056
rect 22468 27004 22520 27056
rect 23112 27004 23164 27056
rect 25412 27047 25464 27056
rect 25412 27013 25421 27047
rect 25421 27013 25455 27047
rect 25455 27013 25464 27047
rect 25412 27004 25464 27013
rect 26792 27004 26844 27056
rect 21456 26979 21508 26988
rect 21456 26945 21465 26979
rect 21465 26945 21499 26979
rect 21499 26945 21508 26979
rect 21456 26936 21508 26945
rect 22652 26979 22704 26988
rect 22652 26945 22661 26979
rect 22661 26945 22695 26979
rect 22695 26945 22704 26979
rect 22652 26936 22704 26945
rect 22928 26979 22980 26988
rect 22928 26945 22937 26979
rect 22937 26945 22971 26979
rect 22971 26945 22980 26979
rect 22928 26936 22980 26945
rect 23020 26979 23072 26988
rect 23020 26945 23029 26979
rect 23029 26945 23063 26979
rect 23063 26945 23072 26979
rect 23020 26936 23072 26945
rect 20628 26843 20680 26852
rect 20628 26809 20637 26843
rect 20637 26809 20671 26843
rect 20671 26809 20680 26843
rect 20628 26800 20680 26809
rect 21824 26843 21876 26852
rect 20168 26775 20220 26784
rect 20168 26741 20177 26775
rect 20177 26741 20211 26775
rect 20211 26741 20220 26775
rect 20168 26732 20220 26741
rect 20444 26732 20496 26784
rect 21824 26809 21833 26843
rect 21833 26809 21867 26843
rect 21867 26809 21876 26843
rect 21824 26800 21876 26809
rect 22284 26800 22336 26852
rect 23664 26936 23716 26988
rect 24400 26936 24452 26988
rect 24676 26936 24728 26988
rect 24768 26936 24820 26988
rect 24952 26936 25004 26988
rect 25136 26936 25188 26988
rect 24492 26911 24544 26920
rect 24492 26877 24501 26911
rect 24501 26877 24535 26911
rect 24535 26877 24544 26911
rect 24492 26868 24544 26877
rect 25228 26868 25280 26920
rect 25872 26979 25924 26988
rect 25872 26945 25881 26979
rect 25881 26945 25915 26979
rect 25915 26945 25924 26979
rect 25872 26936 25924 26945
rect 25964 26936 26016 26988
rect 26240 26936 26292 26988
rect 25596 26800 25648 26852
rect 26148 26843 26200 26852
rect 26148 26809 26157 26843
rect 26157 26809 26191 26843
rect 26191 26809 26200 26843
rect 26148 26800 26200 26809
rect 24216 26775 24268 26784
rect 24216 26741 24225 26775
rect 24225 26741 24259 26775
rect 24259 26741 24268 26775
rect 24216 26732 24268 26741
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 3056 26528 3108 26580
rect 2136 26460 2188 26512
rect 2596 26460 2648 26512
rect 3516 26460 3568 26512
rect 2504 26299 2556 26308
rect 2504 26265 2513 26299
rect 2513 26265 2547 26299
rect 2547 26265 2556 26299
rect 3884 26528 3936 26580
rect 4804 26528 4856 26580
rect 7012 26571 7064 26580
rect 7012 26537 7021 26571
rect 7021 26537 7055 26571
rect 7055 26537 7064 26571
rect 7012 26528 7064 26537
rect 4068 26460 4120 26512
rect 4620 26392 4672 26444
rect 3884 26324 3936 26376
rect 4988 26367 5040 26376
rect 4988 26333 4997 26367
rect 4997 26333 5031 26367
rect 5031 26333 5040 26367
rect 4988 26324 5040 26333
rect 2504 26256 2556 26265
rect 4804 26256 4856 26308
rect 5172 26392 5224 26444
rect 5264 26367 5316 26376
rect 5264 26333 5273 26367
rect 5273 26333 5307 26367
rect 5307 26333 5316 26367
rect 5264 26324 5316 26333
rect 5356 26367 5408 26376
rect 5356 26333 5365 26367
rect 5365 26333 5399 26367
rect 5399 26333 5408 26367
rect 5356 26324 5408 26333
rect 5540 26367 5592 26376
rect 5540 26333 5549 26367
rect 5549 26333 5583 26367
rect 5583 26333 5592 26367
rect 5540 26324 5592 26333
rect 5816 26367 5868 26376
rect 5816 26333 5825 26367
rect 5825 26333 5859 26367
rect 5859 26333 5868 26367
rect 5816 26324 5868 26333
rect 6552 26460 6604 26512
rect 6644 26460 6696 26512
rect 6644 26367 6696 26376
rect 6644 26333 6653 26367
rect 6653 26333 6687 26367
rect 6687 26333 6696 26367
rect 6644 26324 6696 26333
rect 6920 26392 6972 26444
rect 1768 26188 1820 26240
rect 2780 26188 2832 26240
rect 5172 26231 5224 26240
rect 5172 26197 5174 26231
rect 5174 26197 5208 26231
rect 5208 26197 5224 26231
rect 5172 26188 5224 26197
rect 6276 26256 6328 26308
rect 9864 26528 9916 26580
rect 9956 26528 10008 26580
rect 11152 26528 11204 26580
rect 12256 26528 12308 26580
rect 12532 26528 12584 26580
rect 18328 26528 18380 26580
rect 20168 26528 20220 26580
rect 22652 26528 22704 26580
rect 7656 26367 7708 26376
rect 7656 26333 7665 26367
rect 7665 26333 7699 26367
rect 7699 26333 7708 26367
rect 7656 26324 7708 26333
rect 8576 26367 8628 26376
rect 8576 26333 8585 26367
rect 8585 26333 8619 26367
rect 8619 26333 8628 26367
rect 8576 26324 8628 26333
rect 8760 26367 8812 26376
rect 8760 26333 8769 26367
rect 8769 26333 8803 26367
rect 8803 26333 8812 26367
rect 8760 26324 8812 26333
rect 10232 26460 10284 26512
rect 9772 26367 9824 26376
rect 9772 26333 9781 26367
rect 9781 26333 9815 26367
rect 9815 26333 9824 26367
rect 9772 26324 9824 26333
rect 10232 26324 10284 26376
rect 10508 26367 10560 26376
rect 10508 26333 10517 26367
rect 10517 26333 10551 26367
rect 10551 26333 10560 26367
rect 10508 26324 10560 26333
rect 11704 26460 11756 26512
rect 11888 26392 11940 26444
rect 10692 26324 10744 26376
rect 11520 26324 11572 26376
rect 12164 26324 12216 26376
rect 12256 26367 12308 26376
rect 12256 26333 12265 26367
rect 12265 26333 12299 26367
rect 12299 26333 12308 26367
rect 12256 26324 12308 26333
rect 12716 26324 12768 26376
rect 12808 26367 12860 26376
rect 12808 26333 12817 26367
rect 12817 26333 12851 26367
rect 12851 26333 12860 26367
rect 12808 26324 12860 26333
rect 13084 26367 13136 26376
rect 13084 26333 13093 26367
rect 13093 26333 13127 26367
rect 13127 26333 13136 26367
rect 13084 26324 13136 26333
rect 21456 26460 21508 26512
rect 24216 26528 24268 26580
rect 24860 26528 24912 26580
rect 19616 26392 19668 26444
rect 20628 26392 20680 26444
rect 24952 26460 25004 26512
rect 26240 26528 26292 26580
rect 26792 26528 26844 26580
rect 27712 26503 27764 26512
rect 27712 26469 27721 26503
rect 27721 26469 27755 26503
rect 27755 26469 27764 26503
rect 27712 26460 27764 26469
rect 12072 26299 12124 26308
rect 12072 26265 12081 26299
rect 12081 26265 12115 26299
rect 12115 26265 12124 26299
rect 12072 26256 12124 26265
rect 19984 26367 20036 26376
rect 19984 26333 19993 26367
rect 19993 26333 20027 26367
rect 20027 26333 20036 26367
rect 19984 26324 20036 26333
rect 20168 26324 20220 26376
rect 20352 26324 20404 26376
rect 20812 26324 20864 26376
rect 21824 26324 21876 26376
rect 24216 26324 24268 26376
rect 24860 26367 24912 26376
rect 24860 26333 24869 26367
rect 24869 26333 24903 26367
rect 24903 26333 24912 26367
rect 24860 26324 24912 26333
rect 25320 26324 25372 26376
rect 25412 26324 25464 26376
rect 25780 26324 25832 26376
rect 20628 26256 20680 26308
rect 22468 26256 22520 26308
rect 23020 26256 23072 26308
rect 23664 26256 23716 26308
rect 24676 26256 24728 26308
rect 26700 26367 26752 26376
rect 26700 26333 26709 26367
rect 26709 26333 26743 26367
rect 26743 26333 26752 26367
rect 26700 26324 26752 26333
rect 27528 26367 27580 26376
rect 27528 26333 27537 26367
rect 27537 26333 27571 26367
rect 27571 26333 27580 26367
rect 27528 26324 27580 26333
rect 26240 26256 26292 26308
rect 26332 26299 26384 26308
rect 26332 26265 26341 26299
rect 26341 26265 26375 26299
rect 26375 26265 26384 26299
rect 26332 26256 26384 26265
rect 6552 26231 6604 26240
rect 6552 26197 6561 26231
rect 6561 26197 6595 26231
rect 6595 26197 6604 26231
rect 6552 26188 6604 26197
rect 7656 26231 7708 26240
rect 7656 26197 7665 26231
rect 7665 26197 7699 26231
rect 7699 26197 7708 26231
rect 7656 26188 7708 26197
rect 8668 26231 8720 26240
rect 8668 26197 8677 26231
rect 8677 26197 8711 26231
rect 8711 26197 8720 26231
rect 8668 26188 8720 26197
rect 9404 26231 9456 26240
rect 9404 26197 9413 26231
rect 9413 26197 9447 26231
rect 9447 26197 9456 26231
rect 9404 26188 9456 26197
rect 10048 26231 10100 26240
rect 10048 26197 10057 26231
rect 10057 26197 10091 26231
rect 10091 26197 10100 26231
rect 10048 26188 10100 26197
rect 10416 26188 10468 26240
rect 10508 26188 10560 26240
rect 12348 26188 12400 26240
rect 12532 26188 12584 26240
rect 12992 26231 13044 26240
rect 12992 26197 13001 26231
rect 13001 26197 13035 26231
rect 13035 26197 13044 26231
rect 12992 26188 13044 26197
rect 13176 26231 13228 26240
rect 13176 26197 13185 26231
rect 13185 26197 13219 26231
rect 13219 26197 13228 26231
rect 13176 26188 13228 26197
rect 20812 26188 20864 26240
rect 24584 26188 24636 26240
rect 25136 26188 25188 26240
rect 25780 26231 25832 26240
rect 25780 26197 25789 26231
rect 25789 26197 25823 26231
rect 25823 26197 25832 26231
rect 25780 26188 25832 26197
rect 4874 26086 4926 26138
rect 4938 26086 4990 26138
rect 5002 26086 5054 26138
rect 5066 26086 5118 26138
rect 5130 26086 5182 26138
rect 2780 26027 2832 26036
rect 2780 25993 2789 26027
rect 2789 25993 2823 26027
rect 2823 25993 2832 26027
rect 2780 25984 2832 25993
rect 8576 25984 8628 26036
rect 12716 26027 12768 26036
rect 12716 25993 12725 26027
rect 12725 25993 12759 26027
rect 12759 25993 12768 26027
rect 12716 25984 12768 25993
rect 25780 25984 25832 26036
rect 27528 25984 27580 26036
rect 7656 25916 7708 25968
rect 10048 25916 10100 25968
rect 10324 25916 10376 25968
rect 3424 25848 3476 25900
rect 7932 25891 7984 25900
rect 7932 25857 7941 25891
rect 7941 25857 7975 25891
rect 7975 25857 7984 25891
rect 7932 25848 7984 25857
rect 10416 25891 10468 25900
rect 10416 25857 10425 25891
rect 10425 25857 10459 25891
rect 10459 25857 10468 25891
rect 10416 25848 10468 25857
rect 26240 25959 26292 25968
rect 26240 25925 26249 25959
rect 26249 25925 26283 25959
rect 26283 25925 26292 25959
rect 26240 25916 26292 25925
rect 27160 25916 27212 25968
rect 12532 25891 12584 25900
rect 12532 25857 12541 25891
rect 12541 25857 12575 25891
rect 12575 25857 12584 25891
rect 12532 25848 12584 25857
rect 12716 25891 12768 25900
rect 12716 25857 12725 25891
rect 12725 25857 12759 25891
rect 12759 25857 12768 25891
rect 12716 25848 12768 25857
rect 13176 25848 13228 25900
rect 21824 25848 21876 25900
rect 25780 25848 25832 25900
rect 26332 25848 26384 25900
rect 23756 25712 23808 25764
rect 26976 25712 27028 25764
rect 10508 25687 10560 25696
rect 10508 25653 10517 25687
rect 10517 25653 10551 25687
rect 10551 25653 10560 25687
rect 10508 25644 10560 25653
rect 20076 25644 20128 25696
rect 20444 25644 20496 25696
rect 25504 25644 25556 25696
rect 25872 25644 25924 25696
rect 26424 25687 26476 25696
rect 26424 25653 26433 25687
rect 26433 25653 26467 25687
rect 26467 25653 26476 25687
rect 26424 25644 26476 25653
rect 26700 25644 26752 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 20444 25483 20496 25492
rect 20444 25449 20453 25483
rect 20453 25449 20487 25483
rect 20487 25449 20496 25483
rect 20444 25440 20496 25449
rect 20628 25483 20680 25492
rect 20628 25449 20637 25483
rect 20637 25449 20671 25483
rect 20671 25449 20680 25483
rect 20628 25440 20680 25449
rect 20996 25483 21048 25492
rect 20996 25449 21005 25483
rect 21005 25449 21039 25483
rect 21039 25449 21048 25483
rect 20996 25440 21048 25449
rect 2504 25347 2556 25356
rect 2504 25313 2513 25347
rect 2513 25313 2547 25347
rect 2547 25313 2556 25347
rect 2504 25304 2556 25313
rect 2780 25279 2832 25288
rect 2780 25245 2789 25279
rect 2789 25245 2823 25279
rect 2823 25245 2832 25279
rect 2780 25236 2832 25245
rect 5724 25236 5776 25288
rect 10048 25372 10100 25424
rect 10508 25372 10560 25424
rect 6552 25347 6604 25356
rect 6552 25313 6561 25347
rect 6561 25313 6595 25347
rect 6595 25313 6604 25347
rect 6552 25304 6604 25313
rect 7564 25279 7616 25288
rect 7564 25245 7573 25279
rect 7573 25245 7607 25279
rect 7607 25245 7616 25279
rect 7564 25236 7616 25245
rect 5356 25168 5408 25220
rect 7932 25236 7984 25288
rect 8576 25236 8628 25288
rect 8668 25236 8720 25288
rect 9404 25236 9456 25288
rect 10416 25236 10468 25288
rect 11980 25236 12032 25288
rect 12348 25279 12400 25288
rect 12348 25245 12357 25279
rect 12357 25245 12391 25279
rect 12391 25245 12400 25279
rect 12348 25236 12400 25245
rect 12440 25279 12492 25288
rect 12440 25245 12449 25279
rect 12449 25245 12483 25279
rect 12483 25245 12492 25279
rect 12440 25236 12492 25245
rect 13084 25304 13136 25356
rect 15568 25372 15620 25424
rect 15292 25304 15344 25356
rect 12716 25279 12768 25288
rect 12716 25245 12725 25279
rect 12725 25245 12759 25279
rect 12759 25245 12768 25279
rect 12716 25236 12768 25245
rect 15200 25168 15252 25220
rect 15568 25279 15620 25288
rect 15568 25245 15577 25279
rect 15577 25245 15611 25279
rect 15611 25245 15620 25279
rect 15568 25236 15620 25245
rect 16120 25279 16172 25288
rect 16120 25245 16129 25279
rect 16129 25245 16163 25279
rect 16163 25245 16172 25279
rect 16120 25236 16172 25245
rect 22376 25304 22428 25356
rect 21824 25236 21876 25288
rect 23020 25440 23072 25492
rect 27160 25483 27212 25492
rect 27160 25449 27169 25483
rect 27169 25449 27203 25483
rect 27203 25449 27212 25483
rect 27160 25440 27212 25449
rect 22744 25372 22796 25424
rect 24952 25372 25004 25424
rect 23296 25304 23348 25356
rect 22652 25279 22704 25288
rect 22652 25245 22661 25279
rect 22661 25245 22695 25279
rect 22695 25245 22704 25279
rect 22652 25236 22704 25245
rect 23388 25236 23440 25288
rect 25964 25304 26016 25356
rect 25872 25279 25924 25288
rect 25872 25245 25881 25279
rect 25881 25245 25915 25279
rect 25915 25245 25924 25279
rect 25872 25236 25924 25245
rect 26240 25279 26292 25288
rect 26240 25245 26249 25279
rect 26249 25245 26283 25279
rect 26283 25245 26292 25279
rect 26240 25236 26292 25245
rect 16672 25168 16724 25220
rect 20812 25211 20864 25220
rect 20812 25177 20821 25211
rect 20821 25177 20855 25211
rect 20855 25177 20864 25211
rect 20812 25168 20864 25177
rect 22192 25168 22244 25220
rect 23020 25168 23072 25220
rect 3516 25100 3568 25152
rect 7288 25100 7340 25152
rect 7380 25143 7432 25152
rect 7380 25109 7389 25143
rect 7389 25109 7423 25143
rect 7423 25109 7432 25143
rect 7380 25100 7432 25109
rect 8392 25100 8444 25152
rect 9496 25143 9548 25152
rect 9496 25109 9505 25143
rect 9505 25109 9539 25143
rect 9539 25109 9548 25143
rect 9496 25100 9548 25109
rect 10508 25100 10560 25152
rect 12900 25143 12952 25152
rect 12900 25109 12909 25143
rect 12909 25109 12943 25143
rect 12943 25109 12952 25143
rect 12900 25100 12952 25109
rect 16764 25100 16816 25152
rect 20996 25100 21048 25152
rect 23572 25168 23624 25220
rect 24768 25168 24820 25220
rect 23664 25100 23716 25152
rect 26424 25168 26476 25220
rect 27160 25168 27212 25220
rect 26516 25100 26568 25152
rect 27712 25143 27764 25152
rect 27712 25109 27721 25143
rect 27721 25109 27755 25143
rect 27755 25109 27764 25143
rect 27712 25100 27764 25109
rect 4874 24998 4926 25050
rect 4938 24998 4990 25050
rect 5002 24998 5054 25050
rect 5066 24998 5118 25050
rect 5130 24998 5182 25050
rect 11980 24896 12032 24948
rect 12164 24896 12216 24948
rect 16672 24896 16724 24948
rect 10048 24871 10100 24880
rect 10048 24837 10057 24871
rect 10057 24837 10091 24871
rect 10091 24837 10100 24871
rect 10048 24828 10100 24837
rect 5356 24760 5408 24812
rect 7380 24760 7432 24812
rect 3608 24692 3660 24744
rect 4620 24692 4672 24744
rect 8116 24803 8168 24812
rect 8116 24769 8125 24803
rect 8125 24769 8159 24803
rect 8159 24769 8168 24803
rect 8116 24760 8168 24769
rect 8392 24803 8444 24812
rect 8392 24769 8401 24803
rect 8401 24769 8435 24803
rect 8435 24769 8444 24803
rect 8392 24760 8444 24769
rect 9496 24760 9548 24812
rect 10324 24803 10376 24812
rect 10324 24769 10333 24803
rect 10333 24769 10367 24803
rect 10367 24769 10376 24803
rect 10324 24760 10376 24769
rect 10508 24803 10560 24812
rect 10508 24769 10517 24803
rect 10517 24769 10551 24803
rect 10551 24769 10560 24803
rect 10508 24760 10560 24769
rect 4804 24624 4856 24676
rect 8116 24624 8168 24676
rect 10416 24692 10468 24744
rect 11796 24803 11848 24812
rect 11796 24769 11805 24803
rect 11805 24769 11839 24803
rect 11839 24769 11848 24803
rect 11796 24760 11848 24769
rect 12072 24760 12124 24812
rect 11980 24692 12032 24744
rect 5172 24556 5224 24608
rect 8576 24599 8628 24608
rect 8576 24565 8585 24599
rect 8585 24565 8619 24599
rect 8619 24565 8628 24599
rect 8576 24556 8628 24565
rect 9404 24556 9456 24608
rect 9956 24556 10008 24608
rect 10324 24556 10376 24608
rect 13084 24828 13136 24880
rect 13360 24828 13412 24880
rect 12348 24667 12400 24676
rect 12348 24633 12357 24667
rect 12357 24633 12391 24667
rect 12391 24633 12400 24667
rect 13176 24803 13228 24812
rect 13176 24769 13185 24803
rect 13185 24769 13219 24803
rect 13219 24769 13228 24803
rect 13176 24760 13228 24769
rect 14096 24760 14148 24812
rect 15200 24760 15252 24812
rect 15292 24803 15344 24812
rect 15292 24769 15301 24803
rect 15301 24769 15335 24803
rect 15335 24769 15344 24803
rect 15292 24760 15344 24769
rect 15568 24803 15620 24812
rect 15568 24769 15577 24803
rect 15577 24769 15611 24803
rect 15611 24769 15620 24803
rect 15568 24760 15620 24769
rect 16304 24803 16356 24812
rect 16304 24769 16313 24803
rect 16313 24769 16347 24803
rect 16347 24769 16356 24803
rect 16304 24760 16356 24769
rect 16580 24760 16632 24812
rect 16672 24803 16724 24812
rect 16672 24769 16681 24803
rect 16681 24769 16715 24803
rect 16715 24769 16724 24803
rect 16672 24760 16724 24769
rect 16764 24803 16816 24812
rect 16764 24769 16773 24803
rect 16773 24769 16807 24803
rect 16807 24769 16816 24803
rect 16764 24760 16816 24769
rect 20628 24760 20680 24812
rect 21732 24760 21784 24812
rect 22652 24828 22704 24880
rect 24952 24828 25004 24880
rect 16120 24692 16172 24744
rect 12348 24624 12400 24633
rect 15568 24624 15620 24676
rect 17500 24692 17552 24744
rect 24768 24760 24820 24812
rect 25872 24760 25924 24812
rect 22192 24735 22244 24744
rect 22192 24701 22201 24735
rect 22201 24701 22235 24735
rect 22235 24701 22244 24735
rect 22192 24692 22244 24701
rect 12440 24599 12492 24608
rect 12440 24565 12449 24599
rect 12449 24565 12483 24599
rect 12483 24565 12492 24599
rect 12440 24556 12492 24565
rect 13084 24556 13136 24608
rect 15752 24556 15804 24608
rect 15936 24556 15988 24608
rect 17316 24556 17368 24608
rect 21916 24624 21968 24676
rect 22008 24667 22060 24676
rect 22008 24633 22017 24667
rect 22017 24633 22051 24667
rect 22051 24633 22060 24667
rect 22008 24624 22060 24633
rect 17776 24556 17828 24608
rect 23848 24692 23900 24744
rect 24860 24692 24912 24744
rect 24952 24692 25004 24744
rect 25136 24692 25188 24744
rect 26792 24828 26844 24880
rect 26056 24735 26108 24744
rect 26056 24701 26065 24735
rect 26065 24701 26099 24735
rect 26099 24701 26108 24735
rect 26976 24803 27028 24812
rect 26976 24769 26985 24803
rect 26985 24769 27019 24803
rect 27019 24769 27028 24803
rect 26976 24760 27028 24769
rect 26056 24692 26108 24701
rect 26516 24735 26568 24744
rect 26516 24701 26525 24735
rect 26525 24701 26559 24735
rect 26559 24701 26568 24735
rect 26516 24692 26568 24701
rect 25596 24599 25648 24608
rect 25596 24565 25605 24599
rect 25605 24565 25639 24599
rect 25639 24565 25648 24599
rect 25596 24556 25648 24565
rect 25872 24556 25924 24608
rect 27160 24556 27212 24608
rect 27712 24599 27764 24608
rect 27712 24565 27721 24599
rect 27721 24565 27755 24599
rect 27755 24565 27764 24599
rect 27712 24556 27764 24565
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 3608 24395 3660 24404
rect 3608 24361 3617 24395
rect 3617 24361 3651 24395
rect 3651 24361 3660 24395
rect 3608 24352 3660 24361
rect 5356 24395 5408 24404
rect 5356 24361 5365 24395
rect 5365 24361 5399 24395
rect 5399 24361 5408 24395
rect 5356 24352 5408 24361
rect 8116 24352 8168 24404
rect 11980 24395 12032 24404
rect 11980 24361 11989 24395
rect 11989 24361 12023 24395
rect 12023 24361 12032 24395
rect 11980 24352 12032 24361
rect 13176 24352 13228 24404
rect 16212 24352 16264 24404
rect 18144 24352 18196 24404
rect 18604 24352 18656 24404
rect 21732 24395 21784 24404
rect 21732 24361 21741 24395
rect 21741 24361 21775 24395
rect 21775 24361 21784 24395
rect 21732 24352 21784 24361
rect 21824 24352 21876 24404
rect 22008 24352 22060 24404
rect 4068 24284 4120 24336
rect 9312 24327 9364 24336
rect 9312 24293 9321 24327
rect 9321 24293 9355 24327
rect 9355 24293 9364 24327
rect 9312 24284 9364 24293
rect 3516 24216 3568 24268
rect 848 24148 900 24200
rect 1768 24191 1820 24200
rect 1768 24157 1777 24191
rect 1777 24157 1811 24191
rect 1811 24157 1820 24191
rect 1768 24148 1820 24157
rect 2596 24148 2648 24200
rect 2504 24123 2556 24132
rect 2504 24089 2513 24123
rect 2513 24089 2547 24123
rect 2547 24089 2556 24123
rect 3056 24191 3108 24200
rect 3056 24157 3065 24191
rect 3065 24157 3099 24191
rect 3099 24157 3108 24191
rect 3056 24148 3108 24157
rect 4804 24216 4856 24268
rect 7472 24216 7524 24268
rect 2504 24080 2556 24089
rect 4712 24148 4764 24200
rect 5172 24191 5224 24200
rect 5172 24157 5181 24191
rect 5181 24157 5215 24191
rect 5215 24157 5224 24191
rect 5172 24148 5224 24157
rect 4436 24080 4488 24132
rect 4896 24080 4948 24132
rect 7288 24148 7340 24200
rect 8576 24148 8628 24200
rect 9404 24191 9456 24200
rect 9404 24157 9437 24191
rect 9437 24157 9456 24191
rect 9404 24148 9456 24157
rect 9496 24191 9548 24200
rect 9496 24157 9505 24191
rect 9505 24157 9539 24191
rect 9539 24157 9548 24191
rect 9496 24148 9548 24157
rect 9772 24191 9824 24200
rect 9772 24157 9781 24191
rect 9781 24157 9815 24191
rect 9815 24157 9824 24191
rect 9772 24148 9824 24157
rect 9864 24148 9916 24200
rect 10416 24191 10468 24200
rect 10416 24157 10425 24191
rect 10425 24157 10459 24191
rect 10459 24157 10468 24191
rect 10416 24148 10468 24157
rect 11796 24123 11848 24132
rect 11796 24089 11805 24123
rect 11805 24089 11839 24123
rect 11839 24089 11848 24123
rect 11796 24080 11848 24089
rect 12072 24080 12124 24132
rect 12348 24148 12400 24200
rect 12716 24148 12768 24200
rect 12992 24191 13044 24200
rect 12992 24157 13001 24191
rect 13001 24157 13035 24191
rect 13035 24157 13044 24191
rect 12992 24148 13044 24157
rect 13360 24191 13412 24200
rect 13360 24157 13369 24191
rect 13369 24157 13403 24191
rect 13403 24157 13412 24191
rect 13360 24148 13412 24157
rect 14096 24191 14148 24200
rect 14096 24157 14105 24191
rect 14105 24157 14139 24191
rect 14139 24157 14148 24191
rect 14096 24148 14148 24157
rect 17316 24284 17368 24336
rect 17960 24284 18012 24336
rect 18144 24259 18196 24268
rect 18144 24225 18153 24259
rect 18153 24225 18187 24259
rect 18187 24225 18196 24259
rect 18144 24216 18196 24225
rect 19064 24216 19116 24268
rect 19248 24259 19300 24268
rect 19248 24225 19257 24259
rect 19257 24225 19291 24259
rect 19291 24225 19300 24259
rect 19248 24216 19300 24225
rect 23296 24352 23348 24404
rect 24952 24352 25004 24404
rect 26332 24395 26384 24404
rect 26332 24361 26341 24395
rect 26341 24361 26375 24395
rect 26375 24361 26384 24395
rect 26332 24352 26384 24361
rect 21916 24259 21968 24268
rect 21916 24225 21925 24259
rect 21925 24225 21959 24259
rect 21959 24225 21968 24259
rect 21916 24216 21968 24225
rect 22560 24216 22612 24268
rect 17224 24148 17276 24200
rect 17592 24148 17644 24200
rect 17684 24191 17736 24200
rect 17684 24157 17693 24191
rect 17693 24157 17727 24191
rect 17727 24157 17736 24191
rect 17684 24148 17736 24157
rect 17776 24191 17828 24200
rect 17776 24157 17785 24191
rect 17785 24157 17819 24191
rect 17819 24157 17828 24191
rect 17776 24148 17828 24157
rect 18604 24148 18656 24200
rect 20628 24148 20680 24200
rect 21548 24191 21600 24200
rect 21548 24157 21557 24191
rect 21557 24157 21591 24191
rect 21591 24157 21600 24191
rect 21548 24148 21600 24157
rect 14556 24080 14608 24132
rect 15568 24123 15620 24132
rect 15568 24089 15577 24123
rect 15577 24089 15611 24123
rect 15611 24089 15620 24123
rect 15568 24080 15620 24089
rect 16948 24080 17000 24132
rect 18972 24080 19024 24132
rect 1584 24055 1636 24064
rect 1584 24021 1593 24055
rect 1593 24021 1627 24055
rect 1627 24021 1636 24055
rect 1584 24012 1636 24021
rect 5264 24012 5316 24064
rect 16212 24012 16264 24064
rect 16488 24012 16540 24064
rect 16580 24012 16632 24064
rect 17132 24055 17184 24064
rect 17132 24021 17141 24055
rect 17141 24021 17175 24055
rect 17175 24021 17184 24055
rect 17132 24012 17184 24021
rect 17868 24055 17920 24064
rect 17868 24021 17877 24055
rect 17877 24021 17911 24055
rect 17911 24021 17920 24055
rect 17868 24012 17920 24021
rect 18052 24012 18104 24064
rect 21824 24012 21876 24064
rect 22192 24123 22244 24132
rect 22192 24089 22201 24123
rect 22201 24089 22235 24123
rect 22235 24089 22244 24123
rect 22192 24080 22244 24089
rect 23480 24080 23532 24132
rect 24124 24080 24176 24132
rect 24952 24259 25004 24268
rect 24952 24225 24961 24259
rect 24961 24225 24995 24259
rect 24995 24225 25004 24259
rect 24952 24216 25004 24225
rect 25504 24216 25556 24268
rect 25872 24284 25924 24336
rect 24308 24148 24360 24200
rect 24676 24191 24728 24200
rect 24676 24157 24685 24191
rect 24685 24157 24719 24191
rect 24719 24157 24728 24191
rect 24676 24148 24728 24157
rect 23664 24055 23716 24064
rect 23664 24021 23673 24055
rect 23673 24021 23707 24055
rect 23707 24021 23716 24055
rect 24768 24080 24820 24132
rect 25688 24191 25740 24200
rect 25688 24157 25697 24191
rect 25697 24157 25731 24191
rect 25731 24157 25740 24191
rect 25688 24148 25740 24157
rect 25872 24191 25924 24200
rect 25872 24157 25879 24191
rect 25879 24157 25924 24191
rect 25872 24148 25924 24157
rect 26148 24148 26200 24200
rect 25320 24080 25372 24132
rect 23664 24012 23716 24021
rect 24584 24055 24636 24064
rect 24584 24021 24593 24055
rect 24593 24021 24627 24055
rect 24627 24021 24636 24055
rect 24584 24012 24636 24021
rect 25504 24123 25556 24132
rect 25504 24089 25513 24123
rect 25513 24089 25547 24123
rect 25547 24089 25556 24123
rect 25504 24080 25556 24089
rect 25596 24080 25648 24132
rect 26056 24123 26108 24132
rect 26056 24089 26065 24123
rect 26065 24089 26099 24123
rect 26099 24089 26108 24123
rect 26056 24080 26108 24089
rect 26516 24148 26568 24200
rect 26884 24080 26936 24132
rect 27160 24080 27212 24132
rect 27712 24055 27764 24064
rect 27712 24021 27721 24055
rect 27721 24021 27755 24055
rect 27755 24021 27764 24055
rect 27712 24012 27764 24021
rect 4874 23910 4926 23962
rect 4938 23910 4990 23962
rect 5002 23910 5054 23962
rect 5066 23910 5118 23962
rect 5130 23910 5182 23962
rect 1584 23808 1636 23860
rect 1492 23715 1544 23724
rect 1492 23681 1501 23715
rect 1501 23681 1535 23715
rect 1535 23681 1544 23715
rect 1492 23672 1544 23681
rect 3056 23740 3108 23792
rect 2504 23715 2556 23724
rect 2504 23681 2513 23715
rect 2513 23681 2547 23715
rect 2547 23681 2556 23715
rect 2504 23672 2556 23681
rect 3424 23808 3476 23860
rect 3056 23647 3108 23656
rect 3056 23613 3065 23647
rect 3065 23613 3099 23647
rect 3099 23613 3108 23647
rect 3056 23604 3108 23613
rect 2780 23536 2832 23588
rect 3424 23536 3476 23588
rect 4620 23672 4672 23724
rect 4712 23672 4764 23724
rect 5356 23740 5408 23792
rect 4436 23647 4488 23656
rect 4436 23613 4445 23647
rect 4445 23613 4479 23647
rect 4479 23613 4488 23647
rect 4436 23604 4488 23613
rect 4804 23604 4856 23656
rect 8576 23740 8628 23792
rect 10416 23808 10468 23860
rect 8852 23715 8904 23724
rect 8852 23681 8861 23715
rect 8861 23681 8895 23715
rect 8895 23681 8904 23715
rect 8852 23672 8904 23681
rect 9772 23740 9824 23792
rect 9404 23672 9456 23724
rect 12440 23808 12492 23860
rect 16396 23808 16448 23860
rect 17316 23808 17368 23860
rect 17868 23808 17920 23860
rect 18972 23851 19024 23860
rect 18972 23817 18981 23851
rect 18981 23817 19015 23851
rect 19015 23817 19024 23851
rect 18972 23808 19024 23817
rect 21548 23808 21600 23860
rect 24952 23808 25004 23860
rect 25872 23808 25924 23860
rect 26884 23808 26936 23860
rect 12256 23715 12308 23724
rect 12256 23681 12265 23715
rect 12265 23681 12299 23715
rect 12299 23681 12308 23715
rect 12256 23672 12308 23681
rect 12440 23715 12492 23724
rect 12440 23681 12449 23715
rect 12449 23681 12483 23715
rect 12483 23681 12492 23715
rect 12440 23672 12492 23681
rect 13360 23740 13412 23792
rect 14556 23672 14608 23724
rect 15752 23715 15804 23724
rect 15752 23681 15761 23715
rect 15761 23681 15795 23715
rect 15795 23681 15804 23715
rect 15752 23672 15804 23681
rect 15936 23715 15988 23724
rect 15936 23681 15945 23715
rect 15945 23681 15979 23715
rect 15979 23681 15988 23715
rect 15936 23672 15988 23681
rect 16580 23672 16632 23724
rect 17408 23740 17460 23792
rect 22008 23740 22060 23792
rect 23480 23740 23532 23792
rect 25136 23740 25188 23792
rect 25320 23740 25372 23792
rect 10324 23536 10376 23588
rect 12164 23604 12216 23656
rect 17500 23672 17552 23724
rect 17868 23672 17920 23724
rect 18604 23715 18656 23724
rect 18604 23681 18613 23715
rect 18613 23681 18647 23715
rect 18647 23681 18656 23715
rect 18604 23672 18656 23681
rect 18880 23715 18932 23724
rect 18880 23681 18889 23715
rect 18889 23681 18923 23715
rect 18923 23681 18932 23715
rect 18880 23672 18932 23681
rect 19432 23715 19484 23724
rect 19432 23681 19441 23715
rect 19441 23681 19475 23715
rect 19475 23681 19484 23715
rect 19432 23672 19484 23681
rect 19616 23715 19668 23724
rect 19616 23681 19625 23715
rect 19625 23681 19659 23715
rect 19659 23681 19668 23715
rect 19616 23672 19668 23681
rect 20444 23672 20496 23724
rect 21732 23672 21784 23724
rect 17224 23604 17276 23656
rect 17684 23536 17736 23588
rect 2044 23468 2096 23520
rect 5632 23511 5684 23520
rect 5632 23477 5641 23511
rect 5641 23477 5675 23511
rect 5675 23477 5684 23511
rect 5632 23468 5684 23477
rect 12164 23511 12216 23520
rect 12164 23477 12173 23511
rect 12173 23477 12207 23511
rect 12207 23477 12216 23511
rect 12164 23468 12216 23477
rect 12992 23511 13044 23520
rect 12992 23477 13001 23511
rect 13001 23477 13035 23511
rect 13035 23477 13044 23511
rect 12992 23468 13044 23477
rect 15384 23468 15436 23520
rect 15936 23468 15988 23520
rect 16304 23468 16356 23520
rect 16396 23511 16448 23520
rect 16396 23477 16405 23511
rect 16405 23477 16439 23511
rect 16439 23477 16448 23511
rect 16396 23468 16448 23477
rect 16488 23468 16540 23520
rect 17500 23468 17552 23520
rect 17592 23468 17644 23520
rect 18512 23536 18564 23588
rect 17960 23511 18012 23520
rect 17960 23477 17969 23511
rect 17969 23477 18003 23511
rect 18003 23477 18012 23511
rect 17960 23468 18012 23477
rect 18052 23468 18104 23520
rect 23388 23672 23440 23724
rect 23112 23604 23164 23656
rect 24032 23672 24084 23724
rect 25596 23672 25648 23724
rect 25044 23647 25096 23656
rect 25044 23613 25053 23647
rect 25053 23613 25087 23647
rect 25087 23613 25096 23647
rect 25044 23604 25096 23613
rect 25504 23604 25556 23656
rect 23572 23579 23624 23588
rect 23572 23545 23581 23579
rect 23581 23545 23615 23579
rect 23615 23545 23624 23579
rect 27528 23715 27580 23724
rect 27528 23681 27537 23715
rect 27537 23681 27571 23715
rect 27571 23681 27580 23715
rect 27528 23672 27580 23681
rect 23572 23536 23624 23545
rect 23480 23468 23532 23520
rect 24216 23468 24268 23520
rect 27712 23511 27764 23520
rect 27712 23477 27721 23511
rect 27721 23477 27755 23511
rect 27755 23477 27764 23511
rect 27712 23468 27764 23477
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 4620 23264 4672 23316
rect 11796 23264 11848 23316
rect 12992 23307 13044 23316
rect 12992 23273 13001 23307
rect 13001 23273 13035 23307
rect 13035 23273 13044 23307
rect 12992 23264 13044 23273
rect 19616 23307 19668 23316
rect 19616 23273 19625 23307
rect 19625 23273 19659 23307
rect 19659 23273 19668 23307
rect 19616 23264 19668 23273
rect 22192 23264 22244 23316
rect 23388 23264 23440 23316
rect 27528 23264 27580 23316
rect 8852 23196 8904 23248
rect 9312 23196 9364 23248
rect 4620 23060 4672 23112
rect 4712 23060 4764 23112
rect 5264 23128 5316 23180
rect 5540 23171 5592 23180
rect 5540 23137 5549 23171
rect 5549 23137 5583 23171
rect 5583 23137 5592 23171
rect 5540 23128 5592 23137
rect 7288 23128 7340 23180
rect 10324 23128 10376 23180
rect 5448 23060 5500 23112
rect 5632 23103 5684 23112
rect 5632 23069 5641 23103
rect 5641 23069 5675 23103
rect 5675 23069 5684 23103
rect 5632 23060 5684 23069
rect 6184 23103 6236 23112
rect 6184 23069 6193 23103
rect 6193 23069 6227 23103
rect 6227 23069 6236 23103
rect 6184 23060 6236 23069
rect 6276 23060 6328 23112
rect 7472 23103 7524 23112
rect 7472 23069 7481 23103
rect 7481 23069 7515 23103
rect 7515 23069 7524 23103
rect 7472 23060 7524 23069
rect 7932 23103 7984 23112
rect 7932 23069 7941 23103
rect 7941 23069 7975 23103
rect 7975 23069 7984 23103
rect 7932 23060 7984 23069
rect 8852 23060 8904 23112
rect 9312 23060 9364 23112
rect 9496 23060 9548 23112
rect 7288 22992 7340 23044
rect 9956 23103 10008 23112
rect 9956 23069 9965 23103
rect 9965 23069 9999 23103
rect 9999 23069 10008 23103
rect 9956 23060 10008 23069
rect 10232 23103 10284 23112
rect 10232 23069 10241 23103
rect 10241 23069 10275 23103
rect 10275 23069 10284 23103
rect 10232 23060 10284 23069
rect 10508 23103 10560 23112
rect 10508 23069 10517 23103
rect 10517 23069 10551 23103
rect 10551 23069 10560 23103
rect 10508 23060 10560 23069
rect 14280 23128 14332 23180
rect 12256 23060 12308 23112
rect 12532 23060 12584 23112
rect 12624 23103 12676 23112
rect 12624 23069 12633 23103
rect 12633 23069 12667 23103
rect 12667 23069 12676 23103
rect 12624 23060 12676 23069
rect 12900 23103 12952 23112
rect 12900 23069 12909 23103
rect 12909 23069 12943 23103
rect 12943 23069 12952 23103
rect 12900 23060 12952 23069
rect 13268 23103 13320 23112
rect 13268 23069 13277 23103
rect 13277 23069 13311 23103
rect 13311 23069 13320 23103
rect 13268 23060 13320 23069
rect 13544 23060 13596 23112
rect 19340 23196 19392 23248
rect 19432 23196 19484 23248
rect 23664 23196 23716 23248
rect 26240 23196 26292 23248
rect 23480 23128 23532 23180
rect 24400 23171 24452 23180
rect 24400 23137 24409 23171
rect 24409 23137 24443 23171
rect 24443 23137 24452 23171
rect 24400 23128 24452 23137
rect 4620 22924 4672 22976
rect 4896 22924 4948 22976
rect 7840 22967 7892 22976
rect 7840 22933 7849 22967
rect 7849 22933 7883 22967
rect 7883 22933 7892 22967
rect 7840 22924 7892 22933
rect 8024 22967 8076 22976
rect 8024 22933 8033 22967
rect 8033 22933 8067 22967
rect 8067 22933 8076 22967
rect 8024 22924 8076 22933
rect 9772 22924 9824 22976
rect 14096 22924 14148 22976
rect 18696 22967 18748 22976
rect 18696 22933 18705 22967
rect 18705 22933 18739 22967
rect 18739 22933 18748 22967
rect 18696 22924 18748 22933
rect 20352 23103 20404 23112
rect 20352 23069 20361 23103
rect 20361 23069 20395 23103
rect 20395 23069 20404 23103
rect 20352 23060 20404 23069
rect 20444 23103 20496 23112
rect 20444 23069 20453 23103
rect 20453 23069 20487 23103
rect 20487 23069 20496 23103
rect 20444 23060 20496 23069
rect 20812 23060 20864 23112
rect 22744 23060 22796 23112
rect 23848 23060 23900 23112
rect 24032 23103 24084 23112
rect 24032 23069 24041 23103
rect 24041 23069 24075 23103
rect 24075 23069 24084 23103
rect 24032 23060 24084 23069
rect 24216 23103 24268 23112
rect 24216 23069 24225 23103
rect 24225 23069 24259 23103
rect 24259 23069 24268 23103
rect 24216 23060 24268 23069
rect 26148 23060 26200 23112
rect 19340 22992 19392 23044
rect 19432 22967 19484 22976
rect 19432 22933 19441 22967
rect 19441 22933 19475 22967
rect 19475 22933 19484 22967
rect 19432 22924 19484 22933
rect 22468 22992 22520 23044
rect 25136 22992 25188 23044
rect 26884 23035 26936 23044
rect 26884 23001 26893 23035
rect 26893 23001 26927 23035
rect 26927 23001 26936 23035
rect 26884 22992 26936 23001
rect 25504 22924 25556 22976
rect 25964 22924 26016 22976
rect 4874 22822 4926 22874
rect 4938 22822 4990 22874
rect 5002 22822 5054 22874
rect 5066 22822 5118 22874
rect 5130 22822 5182 22874
rect 848 22652 900 22704
rect 2228 22627 2280 22636
rect 2228 22593 2237 22627
rect 2237 22593 2271 22627
rect 2271 22593 2280 22627
rect 2228 22584 2280 22593
rect 3148 22720 3200 22772
rect 7840 22720 7892 22772
rect 3056 22584 3108 22636
rect 8852 22695 8904 22704
rect 8852 22661 8861 22695
rect 8861 22661 8895 22695
rect 8895 22661 8904 22695
rect 8852 22652 8904 22661
rect 9404 22652 9456 22704
rect 3608 22559 3660 22568
rect 3608 22525 3617 22559
rect 3617 22525 3651 22559
rect 3651 22525 3660 22559
rect 3608 22516 3660 22525
rect 5540 22627 5592 22636
rect 5540 22593 5549 22627
rect 5549 22593 5583 22627
rect 5583 22593 5592 22627
rect 5540 22584 5592 22593
rect 6184 22584 6236 22636
rect 5632 22559 5684 22568
rect 5632 22525 5641 22559
rect 5641 22525 5675 22559
rect 5675 22525 5684 22559
rect 5632 22516 5684 22525
rect 6276 22516 6328 22568
rect 8024 22584 8076 22636
rect 9220 22584 9272 22636
rect 10232 22720 10284 22772
rect 13544 22720 13596 22772
rect 17316 22720 17368 22772
rect 17868 22720 17920 22772
rect 19432 22720 19484 22772
rect 20812 22763 20864 22772
rect 20812 22729 20821 22763
rect 20821 22729 20855 22763
rect 20855 22729 20864 22763
rect 20812 22720 20864 22729
rect 26424 22763 26476 22772
rect 26424 22729 26433 22763
rect 26433 22729 26467 22763
rect 26467 22729 26476 22763
rect 26424 22720 26476 22729
rect 9864 22652 9916 22704
rect 9772 22627 9824 22636
rect 9772 22593 9781 22627
rect 9781 22593 9815 22627
rect 9815 22593 9824 22627
rect 9772 22584 9824 22593
rect 10048 22627 10100 22636
rect 10048 22593 10057 22627
rect 10057 22593 10091 22627
rect 10091 22593 10100 22627
rect 10048 22584 10100 22593
rect 10508 22652 10560 22704
rect 14096 22695 14148 22704
rect 14096 22661 14105 22695
rect 14105 22661 14139 22695
rect 14139 22661 14148 22695
rect 14096 22652 14148 22661
rect 16580 22652 16632 22704
rect 10324 22627 10376 22636
rect 10324 22593 10333 22627
rect 10333 22593 10367 22627
rect 10367 22593 10376 22627
rect 10324 22584 10376 22593
rect 2136 22380 2188 22432
rect 2412 22380 2464 22432
rect 3240 22380 3292 22432
rect 12716 22448 12768 22500
rect 13360 22584 13412 22636
rect 13084 22516 13136 22568
rect 13728 22516 13780 22568
rect 18604 22584 18656 22636
rect 20444 22652 20496 22704
rect 26884 22652 26936 22704
rect 20996 22627 21048 22636
rect 20996 22593 21005 22627
rect 21005 22593 21039 22627
rect 21039 22593 21048 22627
rect 20996 22584 21048 22593
rect 13268 22448 13320 22500
rect 20536 22516 20588 22568
rect 22284 22584 22336 22636
rect 25688 22627 25740 22636
rect 25688 22593 25697 22627
rect 25697 22593 25731 22627
rect 25731 22593 25740 22627
rect 25688 22584 25740 22593
rect 25964 22584 26016 22636
rect 26148 22584 26200 22636
rect 3884 22423 3936 22432
rect 3884 22389 3893 22423
rect 3893 22389 3927 22423
rect 3927 22389 3936 22423
rect 3884 22380 3936 22389
rect 6368 22380 6420 22432
rect 7380 22380 7432 22432
rect 7932 22423 7984 22432
rect 7932 22389 7941 22423
rect 7941 22389 7975 22423
rect 7975 22389 7984 22423
rect 7932 22380 7984 22389
rect 9312 22380 9364 22432
rect 10048 22380 10100 22432
rect 12624 22380 12676 22432
rect 12808 22380 12860 22432
rect 14280 22423 14332 22432
rect 14280 22389 14289 22423
rect 14289 22389 14323 22423
rect 14323 22389 14332 22423
rect 14280 22380 14332 22389
rect 16120 22380 16172 22432
rect 27712 22491 27764 22500
rect 27712 22457 27721 22491
rect 27721 22457 27755 22491
rect 27755 22457 27764 22491
rect 27712 22448 27764 22457
rect 17224 22423 17276 22432
rect 17224 22389 17233 22423
rect 17233 22389 17267 22423
rect 17267 22389 17276 22423
rect 17224 22380 17276 22389
rect 19616 22423 19668 22432
rect 19616 22389 19625 22423
rect 19625 22389 19659 22423
rect 19659 22389 19668 22423
rect 19616 22380 19668 22389
rect 25412 22380 25464 22432
rect 25964 22423 26016 22432
rect 25964 22389 25973 22423
rect 25973 22389 26007 22423
rect 26007 22389 26016 22423
rect 25964 22380 26016 22389
rect 26240 22380 26292 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 2228 22083 2280 22092
rect 2228 22049 2237 22083
rect 2237 22049 2271 22083
rect 2271 22049 2280 22083
rect 2228 22040 2280 22049
rect 848 21972 900 22024
rect 3148 22176 3200 22228
rect 4160 22108 4212 22160
rect 3884 22083 3936 22092
rect 3884 22049 3893 22083
rect 3893 22049 3927 22083
rect 3927 22049 3936 22083
rect 3884 22040 3936 22049
rect 4712 22176 4764 22228
rect 7380 22219 7432 22228
rect 7380 22185 7389 22219
rect 7389 22185 7423 22219
rect 7423 22185 7432 22219
rect 7380 22176 7432 22185
rect 20996 22176 21048 22228
rect 21548 22176 21600 22228
rect 26240 22176 26292 22228
rect 14280 22040 14332 22092
rect 3240 22015 3292 22024
rect 3240 21981 3249 22015
rect 3249 21981 3283 22015
rect 3283 21981 3292 22015
rect 3240 21972 3292 21981
rect 3700 21972 3752 22024
rect 3608 21904 3660 21956
rect 3976 21904 4028 21956
rect 2780 21836 2832 21888
rect 2872 21879 2924 21888
rect 2872 21845 2881 21879
rect 2881 21845 2915 21879
rect 2915 21845 2924 21879
rect 2872 21836 2924 21845
rect 3424 21836 3476 21888
rect 4712 21972 4764 22024
rect 7288 22015 7340 22024
rect 7288 21981 7297 22015
rect 7297 21981 7331 22015
rect 7331 21981 7340 22015
rect 7288 21972 7340 21981
rect 7380 21972 7432 22024
rect 9220 22015 9272 22024
rect 9220 21981 9229 22015
rect 9229 21981 9263 22015
rect 9263 21981 9272 22015
rect 9220 21972 9272 21981
rect 9404 22015 9456 22024
rect 9404 21981 9413 22015
rect 9413 21981 9447 22015
rect 9447 21981 9456 22015
rect 9404 21972 9456 21981
rect 9772 22015 9824 22024
rect 9772 21981 9781 22015
rect 9781 21981 9815 22015
rect 9815 21981 9824 22015
rect 9772 21972 9824 21981
rect 12348 21972 12400 22024
rect 13360 22015 13412 22024
rect 13360 21981 13369 22015
rect 13369 21981 13403 22015
rect 13403 21981 13412 22015
rect 13360 21972 13412 21981
rect 13728 21972 13780 22024
rect 14464 21972 14516 22024
rect 16212 22108 16264 22160
rect 17040 22040 17092 22092
rect 17224 21972 17276 22024
rect 17316 22015 17368 22024
rect 17316 21981 17325 22015
rect 17325 21981 17359 22015
rect 17359 21981 17368 22015
rect 17316 21972 17368 21981
rect 24676 21972 24728 22024
rect 26148 22108 26200 22160
rect 25780 22040 25832 22092
rect 26424 22040 26476 22092
rect 25320 22015 25372 22024
rect 25320 21981 25329 22015
rect 25329 21981 25363 22015
rect 25363 21981 25372 22015
rect 25320 21972 25372 21981
rect 25688 21972 25740 22024
rect 14280 21904 14332 21956
rect 16304 21947 16356 21956
rect 16304 21913 16313 21947
rect 16313 21913 16347 21947
rect 16347 21913 16356 21947
rect 16304 21904 16356 21913
rect 25504 21947 25556 21956
rect 25504 21913 25513 21947
rect 25513 21913 25547 21947
rect 25547 21913 25556 21947
rect 25504 21904 25556 21913
rect 4620 21836 4672 21888
rect 13544 21836 13596 21888
rect 14372 21836 14424 21888
rect 15200 21879 15252 21888
rect 15200 21845 15209 21879
rect 15209 21845 15243 21879
rect 15243 21845 15252 21879
rect 15200 21836 15252 21845
rect 16120 21836 16172 21888
rect 17132 21836 17184 21888
rect 17684 21836 17736 21888
rect 25044 21836 25096 21888
rect 25596 21879 25648 21888
rect 25596 21845 25605 21879
rect 25605 21845 25639 21879
rect 25639 21845 25648 21879
rect 25596 21836 25648 21845
rect 25780 21879 25832 21888
rect 25780 21845 25807 21879
rect 25807 21845 25832 21879
rect 25780 21836 25832 21845
rect 26056 21904 26108 21956
rect 26976 21836 27028 21888
rect 4874 21734 4926 21786
rect 4938 21734 4990 21786
rect 5002 21734 5054 21786
rect 5066 21734 5118 21786
rect 5130 21734 5182 21786
rect 2228 21632 2280 21684
rect 4712 21632 4764 21684
rect 13084 21632 13136 21684
rect 14464 21675 14516 21684
rect 14464 21641 14473 21675
rect 14473 21641 14507 21675
rect 14507 21641 14516 21675
rect 14464 21632 14516 21641
rect 19708 21632 19760 21684
rect 23296 21632 23348 21684
rect 24952 21632 25004 21684
rect 25964 21632 26016 21684
rect 26148 21632 26200 21684
rect 19984 21564 20036 21616
rect 20352 21564 20404 21616
rect 25412 21564 25464 21616
rect 26240 21564 26292 21616
rect 2688 21496 2740 21548
rect 3792 21539 3844 21548
rect 3792 21505 3801 21539
rect 3801 21505 3835 21539
rect 3835 21505 3844 21539
rect 3792 21496 3844 21505
rect 3976 21539 4028 21548
rect 3976 21505 3985 21539
rect 3985 21505 4019 21539
rect 4019 21505 4028 21539
rect 3976 21496 4028 21505
rect 4620 21539 4672 21548
rect 4620 21505 4629 21539
rect 4629 21505 4663 21539
rect 4663 21505 4672 21539
rect 4620 21496 4672 21505
rect 4988 21496 5040 21548
rect 7380 21539 7432 21548
rect 7380 21505 7389 21539
rect 7389 21505 7423 21539
rect 7423 21505 7432 21539
rect 7380 21496 7432 21505
rect 12348 21496 12400 21548
rect 2504 21471 2556 21480
rect 2504 21437 2513 21471
rect 2513 21437 2547 21471
rect 2547 21437 2556 21471
rect 2504 21428 2556 21437
rect 5724 21428 5776 21480
rect 7288 21471 7340 21480
rect 7288 21437 7297 21471
rect 7297 21437 7331 21471
rect 7331 21437 7340 21471
rect 7288 21428 7340 21437
rect 8116 21471 8168 21480
rect 8116 21437 8125 21471
rect 8125 21437 8159 21471
rect 8159 21437 8168 21471
rect 8116 21428 8168 21437
rect 12900 21496 12952 21548
rect 13084 21539 13136 21548
rect 13084 21505 13093 21539
rect 13093 21505 13127 21539
rect 13127 21505 13136 21539
rect 13084 21496 13136 21505
rect 13176 21539 13228 21548
rect 13176 21505 13185 21539
rect 13185 21505 13219 21539
rect 13219 21505 13228 21539
rect 13176 21496 13228 21505
rect 13636 21537 13688 21548
rect 13636 21503 13645 21537
rect 13645 21503 13679 21537
rect 13679 21503 13688 21537
rect 13636 21496 13688 21503
rect 14096 21496 14148 21548
rect 14280 21539 14332 21548
rect 14280 21505 14289 21539
rect 14289 21505 14323 21539
rect 14323 21505 14332 21539
rect 14280 21496 14332 21505
rect 14924 21539 14976 21548
rect 14924 21505 14933 21539
rect 14933 21505 14967 21539
rect 14967 21505 14976 21539
rect 14924 21496 14976 21505
rect 15108 21539 15160 21548
rect 15108 21505 15117 21539
rect 15117 21505 15151 21539
rect 15151 21505 15160 21539
rect 15108 21496 15160 21505
rect 16120 21539 16172 21548
rect 16120 21505 16129 21539
rect 16129 21505 16163 21539
rect 16163 21505 16172 21539
rect 16120 21496 16172 21505
rect 16304 21539 16356 21548
rect 16304 21505 16313 21539
rect 16313 21505 16347 21539
rect 16347 21505 16356 21539
rect 16304 21496 16356 21505
rect 17132 21539 17184 21548
rect 17132 21505 17141 21539
rect 17141 21505 17175 21539
rect 17175 21505 17184 21539
rect 17132 21496 17184 21505
rect 16212 21471 16264 21480
rect 16212 21437 16221 21471
rect 16221 21437 16255 21471
rect 16255 21437 16264 21471
rect 16212 21428 16264 21437
rect 17408 21428 17460 21480
rect 18052 21539 18104 21548
rect 18052 21505 18061 21539
rect 18061 21505 18095 21539
rect 18095 21505 18104 21539
rect 18052 21496 18104 21505
rect 17868 21428 17920 21480
rect 19064 21496 19116 21548
rect 21088 21496 21140 21548
rect 23112 21539 23164 21548
rect 23112 21505 23121 21539
rect 23121 21505 23155 21539
rect 23155 21505 23164 21539
rect 23112 21496 23164 21505
rect 12532 21360 12584 21412
rect 13084 21360 13136 21412
rect 13176 21360 13228 21412
rect 13728 21360 13780 21412
rect 12992 21292 13044 21344
rect 13636 21292 13688 21344
rect 14372 21360 14424 21412
rect 17224 21403 17276 21412
rect 17224 21369 17233 21403
rect 17233 21369 17267 21403
rect 17267 21369 17276 21403
rect 17224 21360 17276 21369
rect 17776 21360 17828 21412
rect 19432 21428 19484 21480
rect 22192 21428 22244 21480
rect 22928 21428 22980 21480
rect 24952 21539 25004 21548
rect 24952 21505 24961 21539
rect 24961 21505 24995 21539
rect 24995 21505 25004 21539
rect 24952 21496 25004 21505
rect 25136 21428 25188 21480
rect 21180 21360 21232 21412
rect 22744 21360 22796 21412
rect 25320 21360 25372 21412
rect 25688 21496 25740 21548
rect 27160 21539 27212 21548
rect 27160 21505 27169 21539
rect 27169 21505 27203 21539
rect 27203 21505 27212 21539
rect 27160 21496 27212 21505
rect 25596 21428 25648 21480
rect 26148 21403 26200 21412
rect 26148 21369 26157 21403
rect 26157 21369 26191 21403
rect 26191 21369 26200 21403
rect 26148 21360 26200 21369
rect 26976 21403 27028 21412
rect 26976 21369 26985 21403
rect 26985 21369 27019 21403
rect 27019 21369 27028 21403
rect 26976 21360 27028 21369
rect 16028 21292 16080 21344
rect 19524 21292 19576 21344
rect 19800 21335 19852 21344
rect 19800 21301 19809 21335
rect 19809 21301 19843 21335
rect 19843 21301 19852 21335
rect 19800 21292 19852 21301
rect 21364 21292 21416 21344
rect 23020 21292 23072 21344
rect 25136 21292 25188 21344
rect 25780 21292 25832 21344
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 3792 21088 3844 21140
rect 12348 21131 12400 21140
rect 12348 21097 12357 21131
rect 12357 21097 12391 21131
rect 12391 21097 12400 21131
rect 12348 21088 12400 21097
rect 12716 21088 12768 21140
rect 14004 21088 14056 21140
rect 16304 21088 16356 21140
rect 19064 21088 19116 21140
rect 6368 20995 6420 21004
rect 6368 20961 6377 20995
rect 6377 20961 6411 20995
rect 6411 20961 6420 20995
rect 6368 20952 6420 20961
rect 1032 20884 1084 20936
rect 2688 20884 2740 20936
rect 3700 20884 3752 20936
rect 1492 20859 1544 20868
rect 1492 20825 1501 20859
rect 1501 20825 1535 20859
rect 1535 20825 1544 20859
rect 1492 20816 1544 20825
rect 1768 20816 1820 20868
rect 2136 20816 2188 20868
rect 2504 20816 2556 20868
rect 3424 20816 3476 20868
rect 4068 20884 4120 20936
rect 4620 20884 4672 20936
rect 4988 20927 5040 20936
rect 4988 20893 4997 20927
rect 4997 20893 5031 20927
rect 5031 20893 5040 20927
rect 4988 20884 5040 20893
rect 5632 20927 5684 20936
rect 5632 20893 5641 20927
rect 5641 20893 5675 20927
rect 5675 20893 5684 20927
rect 5632 20884 5684 20893
rect 5724 20927 5776 20936
rect 5724 20893 5733 20927
rect 5733 20893 5767 20927
rect 5767 20893 5776 20927
rect 5724 20884 5776 20893
rect 7748 20952 7800 21004
rect 10600 20927 10652 20936
rect 10600 20893 10609 20927
rect 10609 20893 10643 20927
rect 10643 20893 10652 20927
rect 10600 20884 10652 20893
rect 12992 20995 13044 21004
rect 12992 20961 13001 20995
rect 13001 20961 13035 20995
rect 13035 20961 13044 20995
rect 12992 20952 13044 20961
rect 13084 20927 13136 20936
rect 13084 20893 13093 20927
rect 13093 20893 13127 20927
rect 13127 20893 13136 20927
rect 13084 20884 13136 20893
rect 11152 20816 11204 20868
rect 12256 20816 12308 20868
rect 12992 20816 13044 20868
rect 14188 20884 14240 20936
rect 14372 20884 14424 20936
rect 14648 20884 14700 20936
rect 15108 21020 15160 21072
rect 15200 20995 15252 21004
rect 15200 20961 15209 20995
rect 15209 20961 15243 20995
rect 15243 20961 15252 20995
rect 15200 20952 15252 20961
rect 15108 20927 15160 20936
rect 15108 20893 15117 20927
rect 15117 20893 15151 20927
rect 15151 20893 15160 20927
rect 15108 20884 15160 20893
rect 16212 20952 16264 21004
rect 17132 20952 17184 21004
rect 17408 20995 17460 21004
rect 17408 20961 17417 20995
rect 17417 20961 17451 20995
rect 17451 20961 17460 20995
rect 17408 20952 17460 20961
rect 17868 21020 17920 21072
rect 18604 21020 18656 21072
rect 21180 21088 21232 21140
rect 19524 21063 19576 21072
rect 19524 21029 19533 21063
rect 19533 21029 19567 21063
rect 19567 21029 19576 21063
rect 19524 21020 19576 21029
rect 19616 21063 19668 21072
rect 19616 21029 19625 21063
rect 19625 21029 19659 21063
rect 19659 21029 19668 21063
rect 19616 21020 19668 21029
rect 17776 20995 17828 21004
rect 17776 20961 17785 20995
rect 17785 20961 17819 20995
rect 17819 20961 17828 20995
rect 17776 20952 17828 20961
rect 17960 20952 18012 21004
rect 21364 21020 21416 21072
rect 16120 20884 16172 20936
rect 16580 20884 16632 20936
rect 18604 20927 18656 20936
rect 18604 20893 18613 20927
rect 18613 20893 18647 20927
rect 18647 20893 18656 20927
rect 18604 20884 18656 20893
rect 19064 20884 19116 20936
rect 19616 20884 19668 20936
rect 4068 20748 4120 20800
rect 7104 20791 7156 20800
rect 7104 20757 7113 20791
rect 7113 20757 7147 20791
rect 7147 20757 7156 20791
rect 7104 20748 7156 20757
rect 12532 20791 12584 20800
rect 12532 20757 12541 20791
rect 12541 20757 12575 20791
rect 12575 20757 12584 20791
rect 12532 20748 12584 20757
rect 12624 20748 12676 20800
rect 13360 20748 13412 20800
rect 13912 20748 13964 20800
rect 15476 20816 15528 20868
rect 15844 20791 15896 20800
rect 15844 20757 15853 20791
rect 15853 20757 15887 20791
rect 15887 20757 15896 20791
rect 15844 20748 15896 20757
rect 18328 20816 18380 20868
rect 18512 20816 18564 20868
rect 19156 20816 19208 20868
rect 20076 20927 20128 20936
rect 20076 20893 20085 20927
rect 20085 20893 20119 20927
rect 20119 20893 20128 20927
rect 20076 20884 20128 20893
rect 20168 20927 20220 20936
rect 20168 20893 20177 20927
rect 20177 20893 20211 20927
rect 20211 20893 20220 20927
rect 20168 20884 20220 20893
rect 20536 20927 20588 20936
rect 20536 20893 20545 20927
rect 20545 20893 20579 20927
rect 20579 20893 20588 20927
rect 20536 20884 20588 20893
rect 21088 20927 21140 20936
rect 21088 20893 21097 20927
rect 21097 20893 21131 20927
rect 21131 20893 21140 20927
rect 21548 20995 21600 21004
rect 21548 20961 21557 20995
rect 21557 20961 21591 20995
rect 21591 20961 21600 20995
rect 21548 20952 21600 20961
rect 21088 20884 21140 20893
rect 22008 21020 22060 21072
rect 23940 21088 23992 21140
rect 25044 21131 25096 21140
rect 25044 21097 25053 21131
rect 25053 21097 25087 21131
rect 25087 21097 25096 21131
rect 25044 21088 25096 21097
rect 26056 21088 26108 21140
rect 22560 20995 22612 21004
rect 22560 20961 22569 20995
rect 22569 20961 22603 20995
rect 22603 20961 22612 20995
rect 22560 20952 22612 20961
rect 20260 20816 20312 20868
rect 22100 20927 22152 20936
rect 22100 20893 22109 20927
rect 22109 20893 22143 20927
rect 22143 20893 22152 20927
rect 22100 20884 22152 20893
rect 22192 20927 22244 20936
rect 22192 20893 22201 20927
rect 22201 20893 22235 20927
rect 22235 20893 22244 20927
rect 22192 20884 22244 20893
rect 22376 20927 22428 20936
rect 22376 20893 22385 20927
rect 22385 20893 22419 20927
rect 22419 20893 22428 20927
rect 22376 20884 22428 20893
rect 18052 20748 18104 20800
rect 18696 20748 18748 20800
rect 19524 20748 19576 20800
rect 20352 20791 20404 20800
rect 20352 20757 20361 20791
rect 20361 20757 20395 20791
rect 20395 20757 20404 20791
rect 20352 20748 20404 20757
rect 20904 20748 20956 20800
rect 21916 20791 21968 20800
rect 21916 20757 21925 20791
rect 21925 20757 21959 20791
rect 21959 20757 21968 20791
rect 21916 20748 21968 20757
rect 22284 20816 22336 20868
rect 22744 20927 22796 20936
rect 22744 20893 22753 20927
rect 22753 20893 22787 20927
rect 22787 20893 22796 20927
rect 22744 20884 22796 20893
rect 23020 20927 23072 20936
rect 23020 20893 23029 20927
rect 23029 20893 23063 20927
rect 23063 20893 23072 20927
rect 23020 20884 23072 20893
rect 23296 20927 23348 20936
rect 23296 20893 23305 20927
rect 23305 20893 23339 20927
rect 23339 20893 23348 20927
rect 23296 20884 23348 20893
rect 23388 20927 23440 20936
rect 23388 20893 23397 20927
rect 23397 20893 23431 20927
rect 23431 20893 23440 20927
rect 23388 20884 23440 20893
rect 24308 20884 24360 20936
rect 24400 20884 24452 20936
rect 25320 20927 25372 20936
rect 25320 20893 25329 20927
rect 25329 20893 25363 20927
rect 25363 20893 25372 20927
rect 25320 20884 25372 20893
rect 22192 20748 22244 20800
rect 22376 20748 22428 20800
rect 22744 20748 22796 20800
rect 23572 20859 23624 20868
rect 23572 20825 23581 20859
rect 23581 20825 23615 20859
rect 23615 20825 23624 20859
rect 23572 20816 23624 20825
rect 25872 20816 25924 20868
rect 26608 20816 26660 20868
rect 24216 20748 24268 20800
rect 25044 20791 25096 20800
rect 25044 20757 25069 20791
rect 25069 20757 25096 20791
rect 25044 20748 25096 20757
rect 25228 20791 25280 20800
rect 25228 20757 25237 20791
rect 25237 20757 25271 20791
rect 25271 20757 25280 20791
rect 25228 20748 25280 20757
rect 4874 20646 4926 20698
rect 4938 20646 4990 20698
rect 5002 20646 5054 20698
rect 5066 20646 5118 20698
rect 5130 20646 5182 20698
rect 8392 20544 8444 20596
rect 11152 20544 11204 20596
rect 1952 20519 2004 20528
rect 1952 20485 1961 20519
rect 1961 20485 1995 20519
rect 1995 20485 2004 20519
rect 1952 20476 2004 20485
rect 4160 20476 4212 20528
rect 2596 20408 2648 20460
rect 2688 20451 2740 20460
rect 2688 20417 2697 20451
rect 2697 20417 2731 20451
rect 2731 20417 2740 20451
rect 2688 20408 2740 20417
rect 4804 20451 4856 20460
rect 4804 20417 4813 20451
rect 4813 20417 4847 20451
rect 4847 20417 4856 20451
rect 4804 20408 4856 20417
rect 7104 20519 7156 20528
rect 7104 20485 7113 20519
rect 7113 20485 7147 20519
rect 7147 20485 7156 20519
rect 7104 20476 7156 20485
rect 5724 20408 5776 20460
rect 7564 20408 7616 20460
rect 12716 20544 12768 20596
rect 13084 20544 13136 20596
rect 12532 20476 12584 20528
rect 5632 20340 5684 20392
rect 6460 20340 6512 20392
rect 7748 20383 7800 20392
rect 7748 20349 7757 20383
rect 7757 20349 7791 20383
rect 7791 20349 7800 20383
rect 7748 20340 7800 20349
rect 11796 20383 11848 20392
rect 11796 20349 11805 20383
rect 11805 20349 11839 20383
rect 11839 20349 11848 20383
rect 11796 20340 11848 20349
rect 12348 20383 12400 20392
rect 12348 20349 12357 20383
rect 12357 20349 12391 20383
rect 12391 20349 12400 20383
rect 12348 20340 12400 20349
rect 12716 20408 12768 20460
rect 13360 20408 13412 20460
rect 13452 20451 13504 20460
rect 13452 20417 13461 20451
rect 13461 20417 13495 20451
rect 13495 20417 13504 20451
rect 13452 20408 13504 20417
rect 13544 20451 13596 20460
rect 13544 20417 13553 20451
rect 13553 20417 13587 20451
rect 13587 20417 13596 20451
rect 13544 20408 13596 20417
rect 11980 20272 12032 20324
rect 12440 20272 12492 20324
rect 12808 20340 12860 20392
rect 13912 20451 13964 20460
rect 13912 20417 13921 20451
rect 13921 20417 13955 20451
rect 13955 20417 13964 20451
rect 13912 20408 13964 20417
rect 15016 20544 15068 20596
rect 15568 20544 15620 20596
rect 16396 20544 16448 20596
rect 14096 20476 14148 20528
rect 16304 20476 16356 20528
rect 13084 20272 13136 20324
rect 14556 20451 14608 20460
rect 14556 20417 14565 20451
rect 14565 20417 14599 20451
rect 14599 20417 14608 20451
rect 14556 20408 14608 20417
rect 15292 20451 15344 20460
rect 15292 20417 15301 20451
rect 15301 20417 15335 20451
rect 15335 20417 15344 20451
rect 15292 20408 15344 20417
rect 15384 20451 15436 20460
rect 15384 20417 15393 20451
rect 15393 20417 15427 20451
rect 15427 20417 15436 20451
rect 15384 20408 15436 20417
rect 16212 20451 16264 20460
rect 16212 20417 16221 20451
rect 16221 20417 16255 20451
rect 16255 20417 16264 20451
rect 16212 20408 16264 20417
rect 17040 20451 17092 20460
rect 17040 20417 17049 20451
rect 17049 20417 17083 20451
rect 17083 20417 17092 20451
rect 17040 20408 17092 20417
rect 19616 20544 19668 20596
rect 19892 20544 19944 20596
rect 17684 20451 17736 20460
rect 17684 20417 17693 20451
rect 17693 20417 17727 20451
rect 17727 20417 17736 20451
rect 17684 20408 17736 20417
rect 18512 20476 18564 20528
rect 19524 20519 19576 20528
rect 19524 20485 19533 20519
rect 19533 20485 19567 20519
rect 19567 20485 19576 20519
rect 19524 20476 19576 20485
rect 21088 20544 21140 20596
rect 22008 20587 22060 20596
rect 22008 20553 22033 20587
rect 22033 20553 22060 20587
rect 22008 20544 22060 20553
rect 22192 20587 22244 20596
rect 22192 20553 22201 20587
rect 22201 20553 22235 20587
rect 22235 20553 22244 20587
rect 22192 20544 22244 20553
rect 24216 20587 24268 20596
rect 24216 20553 24225 20587
rect 24225 20553 24259 20587
rect 24259 20553 24268 20587
rect 24216 20544 24268 20553
rect 25044 20544 25096 20596
rect 25872 20544 25924 20596
rect 26240 20544 26292 20596
rect 21824 20519 21876 20528
rect 21824 20485 21833 20519
rect 21833 20485 21867 20519
rect 21867 20485 21876 20519
rect 21824 20476 21876 20485
rect 14372 20383 14424 20392
rect 14372 20349 14381 20383
rect 14381 20349 14415 20383
rect 14415 20349 14424 20383
rect 14372 20340 14424 20349
rect 18236 20340 18288 20392
rect 19156 20451 19208 20460
rect 19156 20417 19165 20451
rect 19165 20417 19199 20451
rect 19199 20417 19208 20451
rect 19156 20408 19208 20417
rect 20628 20408 20680 20460
rect 21180 20408 21232 20460
rect 21364 20451 21416 20460
rect 21364 20417 21373 20451
rect 21373 20417 21407 20451
rect 21407 20417 21416 20451
rect 21364 20408 21416 20417
rect 22836 20476 22888 20528
rect 26976 20476 27028 20528
rect 12808 20204 12860 20256
rect 13452 20204 13504 20256
rect 17132 20272 17184 20324
rect 17316 20272 17368 20324
rect 18236 20204 18288 20256
rect 18512 20204 18564 20256
rect 19248 20383 19300 20392
rect 19248 20349 19257 20383
rect 19257 20349 19291 20383
rect 19291 20349 19300 20383
rect 19248 20340 19300 20349
rect 22560 20383 22612 20392
rect 22560 20349 22569 20383
rect 22569 20349 22603 20383
rect 22603 20349 22612 20383
rect 22560 20340 22612 20349
rect 19156 20272 19208 20324
rect 20628 20272 20680 20324
rect 19892 20204 19944 20256
rect 20076 20204 20128 20256
rect 21916 20204 21968 20256
rect 25780 20451 25832 20460
rect 25780 20417 25789 20451
rect 25789 20417 25823 20451
rect 25823 20417 25832 20451
rect 25780 20408 25832 20417
rect 26148 20408 26200 20460
rect 26240 20451 26292 20460
rect 26240 20417 26249 20451
rect 26249 20417 26283 20451
rect 26283 20417 26292 20451
rect 26240 20408 26292 20417
rect 23756 20204 23808 20256
rect 24032 20247 24084 20256
rect 24032 20213 24041 20247
rect 24041 20213 24075 20247
rect 24075 20213 24084 20247
rect 24032 20204 24084 20213
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 4804 20000 4856 20052
rect 12348 20000 12400 20052
rect 14924 20000 14976 20052
rect 15200 20043 15252 20052
rect 15200 20009 15209 20043
rect 15209 20009 15243 20043
rect 15243 20009 15252 20043
rect 15200 20000 15252 20009
rect 15476 20043 15528 20052
rect 15476 20009 15485 20043
rect 15485 20009 15519 20043
rect 15519 20009 15528 20043
rect 15476 20000 15528 20009
rect 16212 20000 16264 20052
rect 18236 20043 18288 20052
rect 18236 20009 18245 20043
rect 18245 20009 18279 20043
rect 18279 20009 18288 20043
rect 18236 20000 18288 20009
rect 22560 20000 22612 20052
rect 23388 20000 23440 20052
rect 1584 19932 1636 19984
rect 9128 19932 9180 19984
rect 13268 19932 13320 19984
rect 7748 19864 7800 19916
rect 10600 19864 10652 19916
rect 11980 19864 12032 19916
rect 12624 19864 12676 19916
rect 12716 19907 12768 19916
rect 12716 19873 12725 19907
rect 12725 19873 12759 19907
rect 12759 19873 12768 19907
rect 12716 19864 12768 19873
rect 13084 19864 13136 19916
rect 14648 19932 14700 19984
rect 848 19796 900 19848
rect 1952 19796 2004 19848
rect 2228 19839 2280 19848
rect 2228 19805 2237 19839
rect 2237 19805 2271 19839
rect 2271 19805 2280 19839
rect 2228 19796 2280 19805
rect 2412 19839 2464 19848
rect 2412 19805 2421 19839
rect 2421 19805 2455 19839
rect 2455 19805 2464 19839
rect 2412 19796 2464 19805
rect 2872 19796 2924 19848
rect 4160 19796 4212 19848
rect 5356 19796 5408 19848
rect 7380 19796 7432 19848
rect 7564 19839 7616 19848
rect 7564 19805 7573 19839
rect 7573 19805 7607 19839
rect 7607 19805 7616 19839
rect 7564 19796 7616 19805
rect 8116 19796 8168 19848
rect 2688 19728 2740 19780
rect 3700 19728 3752 19780
rect 8392 19728 8444 19780
rect 13268 19796 13320 19848
rect 12256 19728 12308 19780
rect 13452 19796 13504 19848
rect 15016 19864 15068 19916
rect 13728 19796 13780 19848
rect 13912 19796 13964 19848
rect 14372 19839 14424 19848
rect 14372 19805 14381 19839
rect 14381 19805 14415 19839
rect 14415 19805 14424 19839
rect 14372 19796 14424 19805
rect 14556 19839 14608 19848
rect 14556 19805 14565 19839
rect 14565 19805 14599 19839
rect 14599 19805 14608 19839
rect 14556 19796 14608 19805
rect 15108 19839 15160 19848
rect 15108 19805 15117 19839
rect 15117 19805 15151 19839
rect 15151 19805 15160 19839
rect 15108 19796 15160 19805
rect 17960 19864 18012 19916
rect 16396 19839 16448 19848
rect 16396 19805 16405 19839
rect 16405 19805 16439 19839
rect 16439 19805 16448 19839
rect 16396 19796 16448 19805
rect 16580 19771 16632 19780
rect 7840 19660 7892 19712
rect 10048 19703 10100 19712
rect 10048 19669 10057 19703
rect 10057 19669 10091 19703
rect 10091 19669 10100 19703
rect 10048 19660 10100 19669
rect 16580 19737 16589 19771
rect 16589 19737 16623 19771
rect 16623 19737 16632 19771
rect 16580 19728 16632 19737
rect 16764 19728 16816 19780
rect 17224 19728 17276 19780
rect 12900 19660 12952 19712
rect 16396 19660 16448 19712
rect 18144 19660 18196 19712
rect 18788 19839 18840 19848
rect 18788 19805 18797 19839
rect 18797 19805 18831 19839
rect 18831 19805 18840 19839
rect 18788 19796 18840 19805
rect 18972 19864 19024 19916
rect 19340 19932 19392 19984
rect 20168 19975 20220 19984
rect 20168 19941 20177 19975
rect 20177 19941 20211 19975
rect 20211 19941 20220 19975
rect 20168 19932 20220 19941
rect 22100 19932 22152 19984
rect 23296 19932 23348 19984
rect 27160 20000 27212 20052
rect 19708 19839 19760 19848
rect 19708 19805 19717 19839
rect 19717 19805 19751 19839
rect 19751 19805 19760 19839
rect 19708 19796 19760 19805
rect 19892 19864 19944 19916
rect 19984 19796 20036 19848
rect 18880 19771 18932 19780
rect 18880 19737 18915 19771
rect 18915 19737 18932 19771
rect 18880 19728 18932 19737
rect 19524 19728 19576 19780
rect 20076 19660 20128 19712
rect 20352 19907 20404 19916
rect 20352 19873 20361 19907
rect 20361 19873 20395 19907
rect 20395 19873 20404 19907
rect 20352 19864 20404 19873
rect 20260 19796 20312 19848
rect 21548 19839 21600 19848
rect 21548 19805 21557 19839
rect 21557 19805 21591 19839
rect 21591 19805 21600 19839
rect 21548 19796 21600 19805
rect 22652 19907 22704 19916
rect 22652 19873 22661 19907
rect 22661 19873 22695 19907
rect 22695 19873 22704 19907
rect 22652 19864 22704 19873
rect 22836 19864 22888 19916
rect 25320 19864 25372 19916
rect 25964 19864 26016 19916
rect 21916 19839 21968 19848
rect 21916 19805 21925 19839
rect 21925 19805 21959 19839
rect 21959 19805 21968 19839
rect 21916 19796 21968 19805
rect 22008 19839 22060 19848
rect 22008 19805 22017 19839
rect 22017 19805 22051 19839
rect 22051 19805 22060 19839
rect 22008 19796 22060 19805
rect 22192 19796 22244 19848
rect 22468 19839 22520 19848
rect 22468 19805 22477 19839
rect 22477 19805 22511 19839
rect 22511 19805 22520 19839
rect 22468 19796 22520 19805
rect 22560 19796 22612 19848
rect 22928 19796 22980 19848
rect 21824 19771 21876 19780
rect 21824 19737 21833 19771
rect 21833 19737 21867 19771
rect 21867 19737 21876 19771
rect 21824 19728 21876 19737
rect 22100 19660 22152 19712
rect 22192 19703 22244 19712
rect 22192 19669 22201 19703
rect 22201 19669 22235 19703
rect 22235 19669 22244 19703
rect 22192 19660 22244 19669
rect 22376 19728 22428 19780
rect 23296 19796 23348 19848
rect 23664 19728 23716 19780
rect 24032 19771 24084 19780
rect 24032 19737 24041 19771
rect 24041 19737 24075 19771
rect 24075 19737 24084 19771
rect 24032 19728 24084 19737
rect 25872 19771 25924 19780
rect 25872 19737 25881 19771
rect 25881 19737 25915 19771
rect 25915 19737 25924 19771
rect 25872 19728 25924 19737
rect 26608 19728 26660 19780
rect 24124 19660 24176 19712
rect 4874 19558 4926 19610
rect 4938 19558 4990 19610
rect 5002 19558 5054 19610
rect 5066 19558 5118 19610
rect 5130 19558 5182 19610
rect 1584 19499 1636 19508
rect 1584 19465 1593 19499
rect 1593 19465 1627 19499
rect 1627 19465 1636 19499
rect 1584 19456 1636 19465
rect 2872 19456 2924 19508
rect 5540 19456 5592 19508
rect 12256 19456 12308 19508
rect 13636 19456 13688 19508
rect 14004 19456 14056 19508
rect 15568 19456 15620 19508
rect 18512 19499 18564 19508
rect 18512 19465 18521 19499
rect 18521 19465 18555 19499
rect 18555 19465 18564 19499
rect 18512 19456 18564 19465
rect 18788 19456 18840 19508
rect 1400 19363 1452 19372
rect 1400 19329 1409 19363
rect 1409 19329 1443 19363
rect 1443 19329 1452 19363
rect 1400 19320 1452 19329
rect 2228 19320 2280 19372
rect 2412 19320 2464 19372
rect 2044 19295 2096 19304
rect 2044 19261 2053 19295
rect 2053 19261 2087 19295
rect 2087 19261 2096 19295
rect 2044 19252 2096 19261
rect 2688 19295 2740 19304
rect 2688 19261 2697 19295
rect 2697 19261 2731 19295
rect 2731 19261 2740 19295
rect 2688 19252 2740 19261
rect 3608 19295 3660 19304
rect 3608 19261 3617 19295
rect 3617 19261 3651 19295
rect 3651 19261 3660 19295
rect 3608 19252 3660 19261
rect 3700 19295 3752 19304
rect 3700 19261 3709 19295
rect 3709 19261 3743 19295
rect 3743 19261 3752 19295
rect 3700 19252 3752 19261
rect 4712 19363 4764 19372
rect 4712 19329 4721 19363
rect 4721 19329 4755 19363
rect 4755 19329 4764 19363
rect 4712 19320 4764 19329
rect 7840 19363 7892 19372
rect 7840 19329 7849 19363
rect 7849 19329 7883 19363
rect 7883 19329 7892 19363
rect 7840 19320 7892 19329
rect 8116 19363 8168 19372
rect 8116 19329 8125 19363
rect 8125 19329 8159 19363
rect 8159 19329 8168 19363
rect 8116 19320 8168 19329
rect 8392 19320 8444 19372
rect 14188 19388 14240 19440
rect 16396 19388 16448 19440
rect 8944 19320 8996 19372
rect 4804 19184 4856 19236
rect 5264 19252 5316 19304
rect 7564 19184 7616 19236
rect 13728 19320 13780 19372
rect 16120 19320 16172 19372
rect 19064 19388 19116 19440
rect 19340 19431 19392 19440
rect 19340 19397 19349 19431
rect 19349 19397 19383 19431
rect 19383 19397 19392 19431
rect 19340 19388 19392 19397
rect 18696 19363 18748 19372
rect 18696 19329 18705 19363
rect 18705 19329 18739 19363
rect 18739 19329 18748 19363
rect 18696 19320 18748 19329
rect 22100 19456 22152 19508
rect 22560 19456 22612 19508
rect 23572 19456 23624 19508
rect 27620 19499 27672 19508
rect 27620 19465 27629 19499
rect 27629 19465 27663 19499
rect 27663 19465 27672 19499
rect 27620 19456 27672 19465
rect 19708 19388 19760 19440
rect 23664 19388 23716 19440
rect 13360 19184 13412 19236
rect 7932 19159 7984 19168
rect 7932 19125 7941 19159
rect 7941 19125 7975 19159
rect 7975 19125 7984 19159
rect 7932 19116 7984 19125
rect 8208 19116 8260 19168
rect 9680 19116 9732 19168
rect 13176 19159 13228 19168
rect 13176 19125 13185 19159
rect 13185 19125 13219 19159
rect 13219 19125 13228 19159
rect 13176 19116 13228 19125
rect 13268 19116 13320 19168
rect 13820 19252 13872 19304
rect 20076 19320 20128 19372
rect 22468 19363 22520 19372
rect 22468 19329 22477 19363
rect 22477 19329 22511 19363
rect 22511 19329 22520 19363
rect 22468 19320 22520 19329
rect 22652 19320 22704 19372
rect 23020 19320 23072 19372
rect 23296 19363 23348 19372
rect 23296 19329 23305 19363
rect 23305 19329 23339 19363
rect 23339 19329 23348 19363
rect 23296 19320 23348 19329
rect 23388 19363 23440 19372
rect 23388 19329 23397 19363
rect 23397 19329 23431 19363
rect 23431 19329 23440 19363
rect 23388 19320 23440 19329
rect 24032 19320 24084 19372
rect 27804 19363 27856 19372
rect 27804 19329 27813 19363
rect 27813 19329 27847 19363
rect 27847 19329 27856 19363
rect 27804 19320 27856 19329
rect 15200 19184 15252 19236
rect 19524 19184 19576 19236
rect 18880 19159 18932 19168
rect 18880 19125 18889 19159
rect 18889 19125 18923 19159
rect 18923 19125 18932 19159
rect 18880 19116 18932 19125
rect 19708 19159 19760 19168
rect 19708 19125 19717 19159
rect 19717 19125 19751 19159
rect 19751 19125 19760 19159
rect 19708 19116 19760 19125
rect 23480 19116 23532 19168
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 9404 18912 9456 18964
rect 2596 18844 2648 18896
rect 3608 18844 3660 18896
rect 10968 18844 11020 18896
rect 15108 18955 15160 18964
rect 15108 18921 15117 18955
rect 15117 18921 15151 18955
rect 15151 18921 15160 18955
rect 15108 18912 15160 18921
rect 15292 18955 15344 18964
rect 15292 18921 15301 18955
rect 15301 18921 15335 18955
rect 15335 18921 15344 18955
rect 15292 18912 15344 18921
rect 15476 18844 15528 18896
rect 17040 18844 17092 18896
rect 19248 18912 19300 18964
rect 27804 18955 27856 18964
rect 27804 18921 27813 18955
rect 27813 18921 27847 18955
rect 27847 18921 27856 18955
rect 27804 18912 27856 18921
rect 4436 18708 4488 18760
rect 4804 18776 4856 18828
rect 4620 18751 4672 18760
rect 4620 18717 4629 18751
rect 4629 18717 4663 18751
rect 4663 18717 4672 18751
rect 4620 18708 4672 18717
rect 5264 18751 5316 18760
rect 5264 18717 5273 18751
rect 5273 18717 5307 18751
rect 5307 18717 5316 18751
rect 5264 18708 5316 18717
rect 5540 18751 5592 18760
rect 5540 18717 5549 18751
rect 5549 18717 5583 18751
rect 5583 18717 5592 18751
rect 5540 18708 5592 18717
rect 7932 18776 7984 18828
rect 6460 18751 6512 18760
rect 6460 18717 6469 18751
rect 6469 18717 6503 18751
rect 6503 18717 6512 18751
rect 6460 18708 6512 18717
rect 8208 18751 8260 18760
rect 8208 18717 8217 18751
rect 8217 18717 8251 18751
rect 8251 18717 8260 18751
rect 8208 18708 8260 18717
rect 8300 18708 8352 18760
rect 8944 18751 8996 18760
rect 8944 18717 8953 18751
rect 8953 18717 8987 18751
rect 8987 18717 8996 18751
rect 8944 18708 8996 18717
rect 13820 18776 13872 18828
rect 9404 18751 9456 18760
rect 9404 18717 9413 18751
rect 9413 18717 9447 18751
rect 9447 18717 9456 18751
rect 9404 18708 9456 18717
rect 6552 18640 6604 18692
rect 7748 18640 7800 18692
rect 8392 18683 8444 18692
rect 8392 18649 8401 18683
rect 8401 18649 8435 18683
rect 8435 18649 8444 18683
rect 8392 18640 8444 18649
rect 9680 18751 9732 18760
rect 9680 18717 9689 18751
rect 9689 18717 9723 18751
rect 9723 18717 9732 18751
rect 9680 18708 9732 18717
rect 10048 18708 10100 18760
rect 12900 18751 12952 18760
rect 12900 18717 12909 18751
rect 12909 18717 12943 18751
rect 12943 18717 12952 18751
rect 12900 18708 12952 18717
rect 13084 18751 13136 18760
rect 13084 18717 13093 18751
rect 13093 18717 13127 18751
rect 13127 18717 13136 18751
rect 13084 18708 13136 18717
rect 3516 18615 3568 18624
rect 3516 18581 3525 18615
rect 3525 18581 3559 18615
rect 3559 18581 3568 18615
rect 3516 18572 3568 18581
rect 8300 18615 8352 18624
rect 8300 18581 8315 18615
rect 8315 18581 8349 18615
rect 8349 18581 8352 18615
rect 8300 18572 8352 18581
rect 9956 18572 10008 18624
rect 12992 18640 13044 18692
rect 14648 18751 14700 18760
rect 14648 18717 14657 18751
rect 14657 18717 14691 18751
rect 14691 18717 14700 18751
rect 14648 18708 14700 18717
rect 14740 18751 14792 18760
rect 14740 18717 14749 18751
rect 14749 18717 14783 18751
rect 14783 18717 14792 18751
rect 14740 18708 14792 18717
rect 15108 18776 15160 18828
rect 17776 18776 17828 18828
rect 22836 18776 22888 18828
rect 15200 18751 15252 18760
rect 15200 18717 15209 18751
rect 15209 18717 15243 18751
rect 15243 18717 15252 18751
rect 15752 18751 15804 18760
rect 15200 18708 15252 18717
rect 15752 18717 15761 18751
rect 15761 18717 15795 18751
rect 15795 18717 15804 18751
rect 15752 18708 15804 18717
rect 15844 18708 15896 18760
rect 18512 18708 18564 18760
rect 26056 18751 26108 18760
rect 26056 18717 26065 18751
rect 26065 18717 26099 18751
rect 26099 18717 26108 18751
rect 26056 18708 26108 18717
rect 10324 18572 10376 18624
rect 13268 18615 13320 18624
rect 13268 18581 13277 18615
rect 13277 18581 13311 18615
rect 13311 18581 13320 18615
rect 13268 18572 13320 18581
rect 13360 18572 13412 18624
rect 19340 18640 19392 18692
rect 25228 18640 25280 18692
rect 16028 18572 16080 18624
rect 24860 18572 24912 18624
rect 25596 18572 25648 18624
rect 26608 18640 26660 18692
rect 4874 18470 4926 18522
rect 4938 18470 4990 18522
rect 5002 18470 5054 18522
rect 5066 18470 5118 18522
rect 5130 18470 5182 18522
rect 7932 18368 7984 18420
rect 12716 18368 12768 18420
rect 13176 18411 13228 18420
rect 13176 18377 13185 18411
rect 13185 18377 13219 18411
rect 13219 18377 13228 18411
rect 13176 18368 13228 18377
rect 3516 18275 3568 18284
rect 3516 18241 3525 18275
rect 3525 18241 3559 18275
rect 3559 18241 3568 18275
rect 3516 18232 3568 18241
rect 3700 18275 3752 18284
rect 3700 18241 3709 18275
rect 3709 18241 3743 18275
rect 3743 18241 3752 18275
rect 3700 18232 3752 18241
rect 4436 18275 4488 18284
rect 4436 18241 4445 18275
rect 4445 18241 4479 18275
rect 4479 18241 4488 18275
rect 4436 18232 4488 18241
rect 4620 18275 4672 18284
rect 4620 18241 4629 18275
rect 4629 18241 4663 18275
rect 4663 18241 4672 18275
rect 4620 18232 4672 18241
rect 5264 18275 5316 18284
rect 5264 18241 5273 18275
rect 5273 18241 5307 18275
rect 5307 18241 5316 18275
rect 5264 18232 5316 18241
rect 6460 18300 6512 18352
rect 6552 18275 6604 18284
rect 6552 18241 6561 18275
rect 6561 18241 6595 18275
rect 6595 18241 6604 18275
rect 6552 18232 6604 18241
rect 7380 18275 7432 18284
rect 7380 18241 7389 18275
rect 7389 18241 7423 18275
rect 7423 18241 7432 18275
rect 7380 18232 7432 18241
rect 7564 18232 7616 18284
rect 3976 18164 4028 18216
rect 5816 18207 5868 18216
rect 5816 18173 5825 18207
rect 5825 18173 5859 18207
rect 5859 18173 5868 18207
rect 5816 18164 5868 18173
rect 7748 18164 7800 18216
rect 7840 18164 7892 18216
rect 9404 18300 9456 18352
rect 18788 18368 18840 18420
rect 22468 18368 22520 18420
rect 22744 18368 22796 18420
rect 25136 18368 25188 18420
rect 9588 18232 9640 18284
rect 10048 18232 10100 18284
rect 11060 18232 11112 18284
rect 12440 18232 12492 18284
rect 13176 18232 13228 18284
rect 13268 18275 13320 18284
rect 13268 18241 13277 18275
rect 13277 18241 13311 18275
rect 13311 18241 13320 18275
rect 13268 18232 13320 18241
rect 15384 18300 15436 18352
rect 4620 18096 4672 18148
rect 8668 18096 8720 18148
rect 9404 18207 9456 18216
rect 9404 18173 9413 18207
rect 9413 18173 9447 18207
rect 9447 18173 9456 18207
rect 9404 18164 9456 18173
rect 12072 18164 12124 18216
rect 12624 18164 12676 18216
rect 12992 18164 13044 18216
rect 15292 18275 15344 18284
rect 15292 18241 15301 18275
rect 15301 18241 15335 18275
rect 15335 18241 15344 18275
rect 15292 18232 15344 18241
rect 9496 18096 9548 18148
rect 11888 18096 11940 18148
rect 12808 18096 12860 18148
rect 15844 18275 15896 18284
rect 15844 18241 15853 18275
rect 15853 18241 15887 18275
rect 15887 18241 15896 18275
rect 15844 18232 15896 18241
rect 23756 18300 23808 18352
rect 16396 18232 16448 18284
rect 17776 18275 17828 18284
rect 17776 18241 17785 18275
rect 17785 18241 17819 18275
rect 17819 18241 17828 18275
rect 17776 18232 17828 18241
rect 22836 18275 22888 18284
rect 22836 18241 22845 18275
rect 22845 18241 22879 18275
rect 22879 18241 22888 18275
rect 22836 18232 22888 18241
rect 15476 18207 15528 18216
rect 15476 18173 15485 18207
rect 15485 18173 15519 18207
rect 15519 18173 15528 18207
rect 15476 18164 15528 18173
rect 21916 18164 21968 18216
rect 15660 18096 15712 18148
rect 16028 18096 16080 18148
rect 9864 18028 9916 18080
rect 12624 18071 12676 18080
rect 12624 18037 12633 18071
rect 12633 18037 12667 18071
rect 12667 18037 12676 18071
rect 12624 18028 12676 18037
rect 14740 18028 14792 18080
rect 15016 18028 15068 18080
rect 16488 18071 16540 18080
rect 16488 18037 16497 18071
rect 16497 18037 16531 18071
rect 16531 18037 16540 18071
rect 16488 18028 16540 18037
rect 23756 18028 23808 18080
rect 24860 18028 24912 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 2320 17824 2372 17876
rect 2596 17824 2648 17876
rect 11060 17824 11112 17876
rect 13084 17824 13136 17876
rect 15752 17824 15804 17876
rect 8300 17756 8352 17808
rect 9864 17756 9916 17808
rect 9220 17688 9272 17740
rect 1584 17620 1636 17672
rect 7380 17620 7432 17672
rect 7656 17663 7708 17672
rect 7656 17629 7665 17663
rect 7665 17629 7699 17663
rect 7699 17629 7708 17663
rect 7656 17620 7708 17629
rect 7748 17663 7800 17672
rect 7748 17629 7757 17663
rect 7757 17629 7791 17663
rect 7791 17629 7800 17663
rect 7748 17620 7800 17629
rect 9128 17620 9180 17672
rect 9588 17688 9640 17740
rect 9496 17620 9548 17672
rect 8576 17595 8628 17604
rect 8576 17561 8585 17595
rect 8585 17561 8619 17595
rect 8619 17561 8628 17595
rect 8576 17552 8628 17561
rect 9404 17484 9456 17536
rect 10324 17620 10376 17672
rect 10968 17663 11020 17672
rect 10968 17629 10977 17663
rect 10977 17629 11011 17663
rect 11011 17629 11020 17663
rect 10968 17620 11020 17629
rect 12164 17688 12216 17740
rect 12992 17688 13044 17740
rect 11980 17620 12032 17672
rect 12256 17620 12308 17672
rect 15016 17756 15068 17808
rect 16672 17756 16724 17808
rect 10784 17484 10836 17536
rect 11796 17484 11848 17536
rect 14188 17688 14240 17740
rect 13268 17620 13320 17672
rect 13452 17663 13504 17672
rect 13452 17629 13461 17663
rect 13461 17629 13495 17663
rect 13495 17629 13504 17663
rect 13452 17620 13504 17629
rect 14832 17620 14884 17672
rect 16028 17688 16080 17740
rect 16304 17688 16356 17740
rect 19800 17756 19852 17808
rect 20628 17756 20680 17808
rect 15016 17663 15068 17672
rect 15016 17629 15025 17663
rect 15025 17629 15059 17663
rect 15059 17629 15068 17663
rect 15016 17620 15068 17629
rect 16396 17620 16448 17672
rect 16948 17620 17000 17672
rect 17132 17663 17184 17672
rect 17132 17629 17141 17663
rect 17141 17629 17175 17663
rect 17175 17629 17184 17663
rect 17132 17620 17184 17629
rect 17776 17620 17828 17672
rect 19708 17688 19760 17740
rect 20904 17688 20956 17740
rect 22192 17756 22244 17808
rect 14464 17484 14516 17536
rect 14556 17484 14608 17536
rect 16580 17552 16632 17604
rect 17224 17595 17276 17604
rect 17224 17561 17233 17595
rect 17233 17561 17267 17595
rect 17267 17561 17276 17595
rect 17224 17552 17276 17561
rect 17316 17595 17368 17604
rect 17316 17561 17351 17595
rect 17351 17561 17368 17595
rect 18420 17620 18472 17672
rect 17316 17552 17368 17561
rect 18788 17620 18840 17672
rect 19248 17620 19300 17672
rect 20812 17663 20864 17672
rect 20812 17629 20821 17663
rect 20821 17629 20855 17663
rect 20855 17629 20864 17663
rect 22928 17731 22980 17740
rect 22928 17697 22937 17731
rect 22937 17697 22971 17731
rect 22971 17697 22980 17731
rect 22928 17688 22980 17697
rect 23112 17688 23164 17740
rect 23296 17688 23348 17740
rect 20812 17620 20864 17629
rect 19156 17552 19208 17604
rect 21364 17552 21416 17604
rect 23204 17620 23256 17672
rect 23848 17620 23900 17672
rect 23756 17552 23808 17604
rect 26148 17688 26200 17740
rect 24216 17663 24268 17672
rect 24216 17629 24225 17663
rect 24225 17629 24259 17663
rect 24259 17629 24268 17663
rect 24216 17620 24268 17629
rect 24492 17620 24544 17672
rect 16028 17484 16080 17536
rect 16672 17484 16724 17536
rect 16856 17527 16908 17536
rect 16856 17493 16865 17527
rect 16865 17493 16899 17527
rect 16899 17493 16908 17527
rect 16856 17484 16908 17493
rect 17868 17484 17920 17536
rect 17960 17527 18012 17536
rect 17960 17493 17969 17527
rect 17969 17493 18003 17527
rect 18003 17493 18012 17527
rect 17960 17484 18012 17493
rect 18604 17484 18656 17536
rect 18788 17527 18840 17536
rect 18788 17493 18797 17527
rect 18797 17493 18831 17527
rect 18831 17493 18840 17527
rect 18788 17484 18840 17493
rect 20260 17527 20312 17536
rect 20260 17493 20269 17527
rect 20269 17493 20303 17527
rect 20303 17493 20312 17527
rect 20260 17484 20312 17493
rect 20720 17484 20772 17536
rect 20996 17484 21048 17536
rect 21548 17484 21600 17536
rect 23204 17484 23256 17536
rect 24400 17484 24452 17536
rect 24860 17552 24912 17604
rect 24768 17484 24820 17536
rect 4874 17382 4926 17434
rect 4938 17382 4990 17434
rect 5002 17382 5054 17434
rect 5066 17382 5118 17434
rect 5130 17382 5182 17434
rect 2044 17212 2096 17264
rect 2504 17212 2556 17264
rect 848 17144 900 17196
rect 2688 17280 2740 17332
rect 3240 17212 3292 17264
rect 10600 17212 10652 17264
rect 15016 17280 15068 17332
rect 16580 17280 16632 17332
rect 17316 17280 17368 17332
rect 18604 17280 18656 17332
rect 20536 17323 20588 17332
rect 20536 17289 20545 17323
rect 20545 17289 20579 17323
rect 20579 17289 20588 17323
rect 20536 17280 20588 17289
rect 21916 17323 21968 17332
rect 21916 17289 21925 17323
rect 21925 17289 21959 17323
rect 21959 17289 21968 17323
rect 21916 17280 21968 17289
rect 24216 17280 24268 17332
rect 2412 17008 2464 17060
rect 3792 17187 3844 17196
rect 3792 17153 3801 17187
rect 3801 17153 3835 17187
rect 3835 17153 3844 17187
rect 3792 17144 3844 17153
rect 3976 17187 4028 17196
rect 3976 17153 3985 17187
rect 3985 17153 4019 17187
rect 4019 17153 4028 17187
rect 3976 17144 4028 17153
rect 7288 17187 7340 17196
rect 7288 17153 7297 17187
rect 7297 17153 7331 17187
rect 7331 17153 7340 17187
rect 7288 17144 7340 17153
rect 8024 17187 8076 17196
rect 8024 17153 8033 17187
rect 8033 17153 8067 17187
rect 8067 17153 8076 17187
rect 8024 17144 8076 17153
rect 8576 17187 8628 17196
rect 8576 17153 8585 17187
rect 8585 17153 8619 17187
rect 8619 17153 8628 17187
rect 8576 17144 8628 17153
rect 9864 17187 9916 17196
rect 9864 17153 9873 17187
rect 9873 17153 9907 17187
rect 9907 17153 9916 17187
rect 9864 17144 9916 17153
rect 9956 17144 10008 17196
rect 10784 17144 10836 17196
rect 11796 17187 11848 17196
rect 11796 17153 11805 17187
rect 11805 17153 11839 17187
rect 11839 17153 11848 17187
rect 11796 17144 11848 17153
rect 11888 17187 11940 17196
rect 11888 17153 11897 17187
rect 11897 17153 11931 17187
rect 11931 17153 11940 17187
rect 11888 17144 11940 17153
rect 11980 17187 12032 17196
rect 11980 17153 11989 17187
rect 11989 17153 12023 17187
rect 12023 17153 12032 17187
rect 11980 17144 12032 17153
rect 5632 17076 5684 17128
rect 6920 17076 6972 17128
rect 10876 17119 10928 17128
rect 10876 17085 10885 17119
rect 10885 17085 10919 17119
rect 10919 17085 10928 17119
rect 10876 17076 10928 17085
rect 12808 17212 12860 17264
rect 14464 17212 14516 17264
rect 13636 17144 13688 17196
rect 14556 17187 14608 17196
rect 14556 17153 14565 17187
rect 14565 17153 14599 17187
rect 14599 17153 14608 17187
rect 14556 17144 14608 17153
rect 14740 17187 14792 17196
rect 14740 17153 14749 17187
rect 14749 17153 14783 17187
rect 14783 17153 14792 17187
rect 14740 17144 14792 17153
rect 17960 17255 18012 17264
rect 17960 17221 17969 17255
rect 17969 17221 18003 17255
rect 18003 17221 18012 17255
rect 17960 17212 18012 17221
rect 15844 17144 15896 17196
rect 16028 17144 16080 17196
rect 16212 17187 16264 17196
rect 16212 17153 16221 17187
rect 16221 17153 16255 17187
rect 16255 17153 16264 17187
rect 16212 17144 16264 17153
rect 16304 17144 16356 17196
rect 16672 17187 16724 17196
rect 16672 17153 16681 17187
rect 16681 17153 16715 17187
rect 16715 17153 16724 17187
rect 16672 17144 16724 17153
rect 16948 17187 17000 17196
rect 16948 17153 16957 17187
rect 16957 17153 16991 17187
rect 16991 17153 17000 17187
rect 16948 17144 17000 17153
rect 17132 17144 17184 17196
rect 17684 17187 17736 17196
rect 17684 17153 17693 17187
rect 17693 17153 17727 17187
rect 17727 17153 17736 17187
rect 17684 17144 17736 17153
rect 19064 17144 19116 17196
rect 13544 17076 13596 17128
rect 13912 17076 13964 17128
rect 8024 17008 8076 17060
rect 2964 16940 3016 16992
rect 3884 16983 3936 16992
rect 3884 16949 3893 16983
rect 3893 16949 3927 16983
rect 3927 16949 3936 16983
rect 3884 16940 3936 16949
rect 9772 16940 9824 16992
rect 12900 16940 12952 16992
rect 13268 16940 13320 16992
rect 13820 16940 13872 16992
rect 14832 16983 14884 16992
rect 14832 16949 14841 16983
rect 14841 16949 14875 16983
rect 14875 16949 14884 16983
rect 14832 16940 14884 16949
rect 15384 16983 15436 16992
rect 15384 16949 15393 16983
rect 15393 16949 15427 16983
rect 15427 16949 15436 16983
rect 15384 16940 15436 16949
rect 15660 16983 15712 16992
rect 15660 16949 15669 16983
rect 15669 16949 15703 16983
rect 15703 16949 15712 16983
rect 15660 16940 15712 16949
rect 16488 16940 16540 16992
rect 17040 17119 17092 17128
rect 17040 17085 17049 17119
rect 17049 17085 17083 17119
rect 17083 17085 17092 17119
rect 17040 17076 17092 17085
rect 17316 17076 17368 17128
rect 20260 17187 20312 17196
rect 20260 17153 20269 17187
rect 20269 17153 20303 17187
rect 20303 17153 20312 17187
rect 20260 17144 20312 17153
rect 20352 17187 20404 17196
rect 20352 17153 20361 17187
rect 20361 17153 20395 17187
rect 20395 17153 20404 17187
rect 20352 17144 20404 17153
rect 20628 17187 20680 17196
rect 20628 17153 20637 17187
rect 20637 17153 20671 17187
rect 20671 17153 20680 17187
rect 20628 17144 20680 17153
rect 20812 17187 20864 17196
rect 20812 17153 20821 17187
rect 20821 17153 20855 17187
rect 20855 17153 20864 17187
rect 20812 17144 20864 17153
rect 20904 17187 20956 17196
rect 20904 17153 20913 17187
rect 20913 17153 20947 17187
rect 20947 17153 20956 17187
rect 20904 17144 20956 17153
rect 20536 17076 20588 17128
rect 21548 17187 21600 17196
rect 21548 17153 21557 17187
rect 21557 17153 21591 17187
rect 21591 17153 21600 17187
rect 21548 17144 21600 17153
rect 21824 17187 21876 17196
rect 21824 17153 21833 17187
rect 21833 17153 21867 17187
rect 21867 17153 21876 17187
rect 21824 17144 21876 17153
rect 22100 17144 22152 17196
rect 23204 17187 23256 17196
rect 23204 17153 23213 17187
rect 23213 17153 23247 17187
rect 23247 17153 23256 17187
rect 23204 17144 23256 17153
rect 24400 17255 24452 17264
rect 24400 17221 24409 17255
rect 24409 17221 24443 17255
rect 24443 17221 24452 17255
rect 24400 17212 24452 17221
rect 23480 17187 23532 17196
rect 23480 17153 23489 17187
rect 23489 17153 23523 17187
rect 23523 17153 23532 17187
rect 23480 17144 23532 17153
rect 23756 17187 23808 17196
rect 23756 17153 23765 17187
rect 23765 17153 23799 17187
rect 23799 17153 23808 17187
rect 23756 17144 23808 17153
rect 23664 17076 23716 17128
rect 23940 17076 23992 17128
rect 24492 17144 24544 17196
rect 24768 17187 24820 17196
rect 24768 17153 24777 17187
rect 24777 17153 24811 17187
rect 24811 17153 24820 17187
rect 24768 17144 24820 17153
rect 22928 17008 22980 17060
rect 19892 16940 19944 16992
rect 20812 16940 20864 16992
rect 21456 16983 21508 16992
rect 21456 16949 21465 16983
rect 21465 16949 21499 16983
rect 21499 16949 21508 16983
rect 21456 16940 21508 16949
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 2412 16779 2464 16788
rect 2412 16745 2421 16779
rect 2421 16745 2455 16779
rect 2455 16745 2464 16779
rect 2412 16736 2464 16745
rect 7840 16736 7892 16788
rect 9404 16736 9456 16788
rect 13452 16779 13504 16788
rect 13452 16745 13461 16779
rect 13461 16745 13495 16779
rect 13495 16745 13504 16779
rect 13452 16736 13504 16745
rect 13636 16736 13688 16788
rect 2044 16532 2096 16584
rect 2320 16600 2372 16652
rect 3148 16643 3200 16652
rect 3148 16609 3157 16643
rect 3157 16609 3191 16643
rect 3191 16609 3200 16643
rect 3148 16600 3200 16609
rect 3240 16643 3292 16652
rect 3240 16609 3249 16643
rect 3249 16609 3283 16643
rect 3283 16609 3292 16643
rect 3240 16600 3292 16609
rect 2504 16575 2556 16584
rect 2504 16541 2513 16575
rect 2513 16541 2547 16575
rect 2547 16541 2556 16575
rect 2504 16532 2556 16541
rect 2964 16575 3016 16584
rect 2964 16541 2973 16575
rect 2973 16541 3007 16575
rect 3007 16541 3016 16575
rect 2964 16532 3016 16541
rect 4620 16668 4672 16720
rect 5356 16668 5408 16720
rect 10876 16668 10928 16720
rect 15844 16668 15896 16720
rect 17500 16736 17552 16788
rect 16396 16668 16448 16720
rect 3792 16600 3844 16652
rect 3976 16532 4028 16584
rect 4528 16532 4580 16584
rect 5816 16532 5868 16584
rect 8024 16575 8076 16584
rect 8024 16541 8033 16575
rect 8033 16541 8067 16575
rect 8067 16541 8076 16575
rect 8024 16532 8076 16541
rect 8484 16532 8536 16584
rect 9036 16532 9088 16584
rect 9772 16600 9824 16652
rect 12624 16600 12676 16652
rect 13360 16600 13412 16652
rect 15384 16600 15436 16652
rect 17316 16668 17368 16720
rect 17868 16736 17920 16788
rect 18788 16736 18840 16788
rect 19800 16736 19852 16788
rect 22100 16736 22152 16788
rect 25504 16736 25556 16788
rect 12164 16532 12216 16584
rect 12256 16575 12308 16584
rect 12256 16541 12265 16575
rect 12265 16541 12299 16575
rect 12299 16541 12308 16575
rect 12256 16532 12308 16541
rect 6920 16464 6972 16516
rect 7564 16464 7616 16516
rect 8300 16464 8352 16516
rect 8944 16464 8996 16516
rect 4620 16396 4672 16448
rect 5632 16396 5684 16448
rect 8484 16396 8536 16448
rect 8760 16439 8812 16448
rect 8760 16405 8769 16439
rect 8769 16405 8803 16439
rect 8803 16405 8812 16439
rect 8760 16396 8812 16405
rect 11152 16396 11204 16448
rect 12900 16575 12952 16584
rect 12900 16541 12909 16575
rect 12909 16541 12943 16575
rect 12943 16541 12952 16575
rect 12900 16532 12952 16541
rect 13268 16575 13320 16584
rect 13268 16541 13277 16575
rect 13277 16541 13311 16575
rect 13311 16541 13320 16575
rect 13268 16532 13320 16541
rect 12808 16396 12860 16448
rect 15476 16464 15528 16516
rect 18604 16668 18656 16720
rect 17776 16600 17828 16652
rect 18052 16575 18104 16584
rect 18052 16541 18061 16575
rect 18061 16541 18095 16575
rect 18095 16541 18104 16575
rect 18052 16532 18104 16541
rect 18696 16575 18748 16584
rect 18696 16541 18705 16575
rect 18705 16541 18739 16575
rect 18739 16541 18748 16575
rect 18696 16532 18748 16541
rect 19524 16668 19576 16720
rect 20444 16668 20496 16720
rect 20996 16668 21048 16720
rect 19248 16600 19300 16652
rect 20536 16643 20588 16652
rect 20536 16609 20545 16643
rect 20545 16609 20579 16643
rect 20579 16609 20588 16643
rect 20536 16600 20588 16609
rect 20720 16643 20772 16652
rect 20720 16609 20729 16643
rect 20729 16609 20763 16643
rect 20763 16609 20772 16643
rect 20720 16600 20772 16609
rect 19064 16532 19116 16584
rect 20444 16575 20496 16584
rect 20444 16541 20453 16575
rect 20453 16541 20487 16575
rect 20487 16541 20496 16575
rect 20444 16532 20496 16541
rect 21456 16600 21508 16652
rect 16028 16396 16080 16448
rect 17224 16439 17276 16448
rect 17224 16405 17233 16439
rect 17233 16405 17267 16439
rect 17267 16405 17276 16439
rect 17224 16396 17276 16405
rect 18052 16439 18104 16448
rect 18052 16405 18061 16439
rect 18061 16405 18095 16439
rect 18095 16405 18104 16439
rect 18052 16396 18104 16405
rect 21088 16464 21140 16516
rect 22100 16575 22152 16584
rect 22100 16541 22109 16575
rect 22109 16541 22143 16575
rect 22143 16541 22152 16575
rect 22100 16532 22152 16541
rect 26148 16643 26200 16652
rect 26148 16609 26157 16643
rect 26157 16609 26191 16643
rect 26191 16609 26200 16643
rect 26148 16600 26200 16609
rect 21640 16464 21692 16516
rect 19708 16396 19760 16448
rect 20996 16396 21048 16448
rect 21272 16396 21324 16448
rect 21364 16439 21416 16448
rect 21364 16405 21373 16439
rect 21373 16405 21407 16439
rect 21407 16405 21416 16439
rect 21364 16396 21416 16405
rect 23388 16439 23440 16448
rect 23388 16405 23397 16439
rect 23397 16405 23431 16439
rect 23431 16405 23440 16439
rect 23388 16396 23440 16405
rect 25320 16464 25372 16516
rect 26608 16507 26660 16516
rect 26608 16473 26617 16507
rect 26617 16473 26651 16507
rect 26651 16473 26660 16507
rect 26608 16464 26660 16473
rect 24860 16396 24912 16448
rect 4874 16294 4926 16346
rect 4938 16294 4990 16346
rect 5002 16294 5054 16346
rect 5066 16294 5118 16346
rect 5130 16294 5182 16346
rect 2504 16056 2556 16108
rect 3884 16099 3936 16108
rect 3884 16065 3893 16099
rect 3893 16065 3927 16099
rect 3927 16065 3936 16099
rect 3884 16056 3936 16065
rect 4620 16099 4672 16108
rect 4620 16065 4629 16099
rect 4629 16065 4663 16099
rect 4663 16065 4672 16099
rect 4620 16056 4672 16065
rect 4896 16099 4948 16108
rect 4896 16065 4905 16099
rect 4905 16065 4939 16099
rect 4939 16065 4948 16099
rect 4896 16056 4948 16065
rect 5356 16099 5408 16108
rect 5356 16065 5365 16099
rect 5365 16065 5399 16099
rect 5399 16065 5408 16099
rect 5356 16056 5408 16065
rect 6920 16192 6972 16244
rect 8760 16124 8812 16176
rect 16672 16192 16724 16244
rect 16948 16192 17000 16244
rect 18512 16192 18564 16244
rect 18788 16192 18840 16244
rect 19064 16192 19116 16244
rect 22008 16192 22060 16244
rect 25320 16235 25372 16244
rect 25320 16201 25329 16235
rect 25329 16201 25363 16235
rect 25363 16201 25372 16235
rect 25320 16192 25372 16201
rect 25688 16192 25740 16244
rect 7288 16056 7340 16108
rect 8208 16056 8260 16108
rect 8944 16056 8996 16108
rect 9036 16099 9088 16108
rect 9036 16065 9045 16099
rect 9045 16065 9079 16099
rect 9079 16065 9088 16099
rect 9036 16056 9088 16065
rect 2228 15988 2280 16040
rect 4528 16031 4580 16040
rect 4528 15997 4537 16031
rect 4537 15997 4571 16031
rect 4571 15997 4580 16031
rect 4528 15988 4580 15997
rect 8852 16031 8904 16040
rect 8852 15997 8861 16031
rect 8861 15997 8895 16031
rect 8895 15997 8904 16031
rect 8852 15988 8904 15997
rect 9772 16099 9824 16108
rect 9772 16065 9781 16099
rect 9781 16065 9815 16099
rect 9815 16065 9824 16099
rect 9772 16056 9824 16065
rect 12808 16167 12860 16176
rect 12808 16133 12817 16167
rect 12817 16133 12851 16167
rect 12851 16133 12860 16167
rect 12808 16124 12860 16133
rect 12992 16124 13044 16176
rect 18236 16124 18288 16176
rect 18696 16124 18748 16176
rect 22192 16124 22244 16176
rect 18052 16056 18104 16108
rect 18512 16099 18564 16108
rect 18512 16065 18521 16099
rect 18521 16065 18555 16099
rect 18555 16065 18564 16099
rect 18512 16056 18564 16065
rect 20536 16099 20588 16108
rect 20536 16065 20545 16099
rect 20545 16065 20579 16099
rect 20579 16065 20588 16099
rect 20536 16056 20588 16065
rect 20812 16099 20864 16108
rect 20812 16065 20821 16099
rect 20821 16065 20855 16099
rect 20855 16065 20864 16099
rect 20812 16056 20864 16065
rect 21272 16099 21324 16108
rect 21272 16065 21281 16099
rect 21281 16065 21315 16099
rect 21315 16065 21324 16099
rect 21272 16056 21324 16065
rect 21640 16056 21692 16108
rect 16856 15988 16908 16040
rect 17960 16031 18012 16040
rect 17960 15997 17969 16031
rect 17969 15997 18003 16031
rect 18003 15997 18012 16031
rect 17960 15988 18012 15997
rect 18328 15988 18380 16040
rect 20996 15988 21048 16040
rect 17040 15920 17092 15972
rect 17408 15920 17460 15972
rect 18696 15920 18748 15972
rect 22560 16056 22612 16108
rect 22744 16099 22796 16108
rect 22744 16065 22753 16099
rect 22753 16065 22787 16099
rect 22787 16065 22796 16099
rect 22744 16056 22796 16065
rect 22928 16099 22980 16108
rect 22928 16065 22937 16099
rect 22937 16065 22971 16099
rect 22971 16065 22980 16099
rect 22928 16056 22980 16065
rect 23388 16124 23440 16176
rect 25504 16124 25556 16176
rect 22100 15988 22152 16040
rect 2320 15852 2372 15904
rect 8300 15852 8352 15904
rect 12808 15895 12860 15904
rect 12808 15861 12817 15895
rect 12817 15861 12851 15895
rect 12851 15861 12860 15895
rect 12808 15852 12860 15861
rect 18144 15895 18196 15904
rect 18144 15861 18153 15895
rect 18153 15861 18187 15895
rect 18187 15861 18196 15895
rect 18144 15852 18196 15861
rect 18604 15852 18656 15904
rect 19340 15852 19392 15904
rect 19800 15852 19852 15904
rect 21088 15852 21140 15904
rect 21364 15852 21416 15904
rect 23572 16099 23624 16108
rect 23572 16065 23581 16099
rect 23581 16065 23615 16099
rect 23615 16065 23624 16099
rect 23572 16056 23624 16065
rect 23388 15988 23440 16040
rect 23848 16056 23900 16108
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 7564 15691 7616 15700
rect 7564 15657 7573 15691
rect 7573 15657 7607 15691
rect 7607 15657 7616 15691
rect 7564 15648 7616 15657
rect 16948 15648 17000 15700
rect 18696 15648 18748 15700
rect 4620 15512 4672 15564
rect 1400 15487 1452 15496
rect 1400 15453 1409 15487
rect 1409 15453 1443 15487
rect 1443 15453 1452 15487
rect 1400 15444 1452 15453
rect 2780 15487 2832 15496
rect 2780 15453 2789 15487
rect 2789 15453 2823 15487
rect 2823 15453 2832 15487
rect 2780 15444 2832 15453
rect 3240 15444 3292 15496
rect 2044 15376 2096 15428
rect 4896 15487 4948 15496
rect 4896 15453 4905 15487
rect 4905 15453 4939 15487
rect 4939 15453 4948 15487
rect 4896 15444 4948 15453
rect 5356 15444 5408 15496
rect 8484 15580 8536 15632
rect 8852 15580 8904 15632
rect 19432 15623 19484 15632
rect 19432 15589 19441 15623
rect 19441 15589 19475 15623
rect 19475 15589 19484 15623
rect 19432 15580 19484 15589
rect 8300 15512 8352 15564
rect 7932 15444 7984 15496
rect 8392 15444 8444 15496
rect 8576 15487 8628 15496
rect 8576 15453 8585 15487
rect 8585 15453 8619 15487
rect 8619 15453 8628 15487
rect 8576 15444 8628 15453
rect 8760 15487 8812 15496
rect 8760 15453 8769 15487
rect 8769 15453 8803 15487
rect 8803 15453 8812 15487
rect 8760 15444 8812 15453
rect 21088 15691 21140 15700
rect 21088 15657 21097 15691
rect 21097 15657 21131 15691
rect 21131 15657 21140 15691
rect 21088 15648 21140 15657
rect 21272 15648 21324 15700
rect 21364 15623 21416 15632
rect 21364 15589 21373 15623
rect 21373 15589 21407 15623
rect 21407 15589 21416 15623
rect 21364 15580 21416 15589
rect 9036 15512 9088 15564
rect 19616 15555 19668 15564
rect 19616 15521 19625 15555
rect 19625 15521 19659 15555
rect 19659 15521 19668 15555
rect 19616 15512 19668 15521
rect 9864 15487 9916 15496
rect 9864 15453 9873 15487
rect 9873 15453 9907 15487
rect 9907 15453 9916 15487
rect 9864 15444 9916 15453
rect 19432 15487 19484 15496
rect 19432 15453 19441 15487
rect 19441 15453 19475 15487
rect 19475 15453 19484 15487
rect 19432 15444 19484 15453
rect 19800 15487 19852 15496
rect 19800 15453 19809 15487
rect 19809 15453 19843 15487
rect 19843 15453 19852 15487
rect 19800 15444 19852 15453
rect 20996 15512 21048 15564
rect 20720 15487 20772 15496
rect 20720 15453 20729 15487
rect 20729 15453 20763 15487
rect 20763 15453 20772 15487
rect 20720 15444 20772 15453
rect 9128 15376 9180 15428
rect 21272 15487 21324 15496
rect 21272 15453 21281 15487
rect 21281 15453 21315 15487
rect 21315 15453 21324 15487
rect 21272 15444 21324 15453
rect 21456 15487 21508 15496
rect 21456 15453 21465 15487
rect 21465 15453 21499 15487
rect 21499 15453 21508 15487
rect 21456 15444 21508 15453
rect 21640 15444 21692 15496
rect 23572 15648 23624 15700
rect 24492 15648 24544 15700
rect 24584 15691 24636 15700
rect 24584 15657 24593 15691
rect 24593 15657 24627 15691
rect 24627 15657 24636 15691
rect 24584 15648 24636 15657
rect 22376 15580 22428 15632
rect 22652 15580 22704 15632
rect 22928 15580 22980 15632
rect 24584 15512 24636 15564
rect 22100 15444 22152 15496
rect 3240 15308 3292 15360
rect 4804 15351 4856 15360
rect 4804 15317 4813 15351
rect 4813 15317 4847 15351
rect 4847 15317 4856 15351
rect 4804 15308 4856 15317
rect 18604 15308 18656 15360
rect 23204 15444 23256 15496
rect 23756 15487 23808 15496
rect 23756 15453 23765 15487
rect 23765 15453 23799 15487
rect 23799 15453 23808 15487
rect 23756 15444 23808 15453
rect 24032 15487 24084 15496
rect 24032 15453 24041 15487
rect 24041 15453 24075 15487
rect 24075 15453 24084 15487
rect 24032 15444 24084 15453
rect 24216 15487 24268 15496
rect 24216 15453 24225 15487
rect 24225 15453 24259 15487
rect 24259 15453 24268 15487
rect 24216 15444 24268 15453
rect 24860 15419 24912 15428
rect 24860 15385 24869 15419
rect 24869 15385 24903 15419
rect 24903 15385 24912 15419
rect 24860 15376 24912 15385
rect 25136 15487 25188 15496
rect 25136 15453 25145 15487
rect 25145 15453 25179 15487
rect 25179 15453 25188 15487
rect 25136 15444 25188 15453
rect 4874 15206 4926 15258
rect 4938 15206 4990 15258
rect 5002 15206 5054 15258
rect 5066 15206 5118 15258
rect 5130 15206 5182 15258
rect 2780 15104 2832 15156
rect 12808 15104 12860 15156
rect 14832 15104 14884 15156
rect 18512 15104 18564 15156
rect 20720 15104 20772 15156
rect 5356 15036 5408 15088
rect 9864 15079 9916 15088
rect 9864 15045 9873 15079
rect 9873 15045 9907 15079
rect 9907 15045 9916 15079
rect 9864 15036 9916 15045
rect 10232 15036 10284 15088
rect 22008 15036 22060 15088
rect 2044 14900 2096 14952
rect 3148 14968 3200 15020
rect 7656 14968 7708 15020
rect 8300 14968 8352 15020
rect 8392 15011 8444 15020
rect 8392 14977 8401 15011
rect 8401 14977 8435 15011
rect 8435 14977 8444 15011
rect 8392 14968 8444 14977
rect 11520 15011 11572 15020
rect 11520 14977 11529 15011
rect 11529 14977 11563 15011
rect 11563 14977 11572 15011
rect 11520 14968 11572 14977
rect 11704 15011 11756 15020
rect 11704 14977 11713 15011
rect 11713 14977 11747 15011
rect 11747 14977 11756 15011
rect 11704 14968 11756 14977
rect 11888 15011 11940 15020
rect 11888 14977 11897 15011
rect 11897 14977 11931 15011
rect 11931 14977 11940 15011
rect 11888 14968 11940 14977
rect 12624 15011 12676 15020
rect 12624 14977 12633 15011
rect 12633 14977 12667 15011
rect 12667 14977 12676 15011
rect 12624 14968 12676 14977
rect 13636 14968 13688 15020
rect 14280 14968 14332 15020
rect 5448 14943 5500 14952
rect 5448 14909 5457 14943
rect 5457 14909 5491 14943
rect 5491 14909 5500 14943
rect 5448 14900 5500 14909
rect 4804 14832 4856 14884
rect 3148 14764 3200 14816
rect 4620 14764 4672 14816
rect 6184 14764 6236 14816
rect 12256 14875 12308 14884
rect 12256 14841 12265 14875
rect 12265 14841 12299 14875
rect 12299 14841 12308 14875
rect 12256 14832 12308 14841
rect 13176 14900 13228 14952
rect 14004 14900 14056 14952
rect 15200 14943 15252 14952
rect 15200 14909 15209 14943
rect 15209 14909 15243 14943
rect 15243 14909 15252 14943
rect 15200 14900 15252 14909
rect 15292 14900 15344 14952
rect 18144 14968 18196 15020
rect 19616 14968 19668 15020
rect 21272 14968 21324 15020
rect 16856 14900 16908 14952
rect 18328 14900 18380 14952
rect 21456 14900 21508 14952
rect 21824 14900 21876 14952
rect 13452 14832 13504 14884
rect 24584 14968 24636 15020
rect 14188 14764 14240 14816
rect 15568 14807 15620 14816
rect 15568 14773 15577 14807
rect 15577 14773 15611 14807
rect 15611 14773 15620 14807
rect 15568 14764 15620 14773
rect 15936 14764 15988 14816
rect 20076 14764 20128 14816
rect 23020 14764 23072 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 11980 14560 12032 14612
rect 4712 14492 4764 14544
rect 8392 14492 8444 14544
rect 12624 14560 12676 14612
rect 14188 14560 14240 14612
rect 15108 14560 15160 14612
rect 4252 14424 4304 14476
rect 5908 14424 5960 14476
rect 11888 14424 11940 14476
rect 12716 14424 12768 14476
rect 2780 14399 2832 14408
rect 2780 14365 2789 14399
rect 2789 14365 2823 14399
rect 2823 14365 2832 14399
rect 2780 14356 2832 14365
rect 3240 14399 3292 14408
rect 3240 14365 3249 14399
rect 3249 14365 3283 14399
rect 3283 14365 3292 14399
rect 3240 14356 3292 14365
rect 3608 14356 3660 14408
rect 4160 14399 4212 14408
rect 4160 14365 4169 14399
rect 4169 14365 4203 14399
rect 4203 14365 4212 14399
rect 4160 14356 4212 14365
rect 4620 14356 4672 14408
rect 4804 14356 4856 14408
rect 5448 14399 5500 14408
rect 5448 14365 5457 14399
rect 5457 14365 5491 14399
rect 5491 14365 5500 14399
rect 5448 14356 5500 14365
rect 6184 14399 6236 14408
rect 6184 14365 6193 14399
rect 6193 14365 6227 14399
rect 6227 14365 6236 14399
rect 6184 14356 6236 14365
rect 6736 14399 6788 14408
rect 6736 14365 6745 14399
rect 6745 14365 6779 14399
rect 6779 14365 6788 14399
rect 6736 14356 6788 14365
rect 11152 14399 11204 14408
rect 11152 14365 11161 14399
rect 11161 14365 11195 14399
rect 11195 14365 11204 14399
rect 11152 14356 11204 14365
rect 11244 14399 11296 14408
rect 11244 14365 11253 14399
rect 11253 14365 11287 14399
rect 11287 14365 11296 14399
rect 11244 14356 11296 14365
rect 13544 14399 13596 14408
rect 13544 14365 13553 14399
rect 13553 14365 13587 14399
rect 13587 14365 13596 14399
rect 13544 14356 13596 14365
rect 13636 14399 13688 14408
rect 13636 14365 13645 14399
rect 13645 14365 13679 14399
rect 13679 14365 13688 14399
rect 13636 14356 13688 14365
rect 15660 14560 15712 14612
rect 17132 14560 17184 14612
rect 24860 14560 24912 14612
rect 25412 14560 25464 14612
rect 23756 14492 23808 14544
rect 24768 14492 24820 14544
rect 17040 14467 17092 14476
rect 17040 14433 17049 14467
rect 17049 14433 17083 14467
rect 17083 14433 17092 14467
rect 17040 14424 17092 14433
rect 17224 14424 17276 14476
rect 19156 14424 19208 14476
rect 20720 14424 20772 14476
rect 22376 14424 22428 14476
rect 25136 14424 25188 14476
rect 2320 14220 2372 14272
rect 3700 14220 3752 14272
rect 12900 14288 12952 14340
rect 12256 14220 12308 14272
rect 12992 14263 13044 14272
rect 12992 14229 13001 14263
rect 13001 14229 13035 14263
rect 13035 14229 13044 14263
rect 12992 14220 13044 14229
rect 14648 14220 14700 14272
rect 14832 14399 14884 14408
rect 14832 14365 14841 14399
rect 14841 14365 14875 14399
rect 14875 14365 14884 14399
rect 14832 14356 14884 14365
rect 15016 14399 15068 14408
rect 15016 14365 15025 14399
rect 15025 14365 15059 14399
rect 15059 14365 15068 14399
rect 15016 14356 15068 14365
rect 15292 14356 15344 14408
rect 15660 14356 15712 14408
rect 16672 14399 16724 14408
rect 16672 14365 16681 14399
rect 16681 14365 16715 14399
rect 16715 14365 16724 14399
rect 16672 14356 16724 14365
rect 16764 14399 16816 14408
rect 16764 14365 16773 14399
rect 16773 14365 16807 14399
rect 16807 14365 16816 14399
rect 16764 14356 16816 14365
rect 17868 14356 17920 14408
rect 18420 14356 18472 14408
rect 19064 14356 19116 14408
rect 15660 14220 15712 14272
rect 18236 14288 18288 14340
rect 19708 14288 19760 14340
rect 20628 14288 20680 14340
rect 24584 14399 24636 14408
rect 24584 14365 24593 14399
rect 24593 14365 24627 14399
rect 24627 14365 24636 14399
rect 24584 14356 24636 14365
rect 27804 14399 27856 14408
rect 27804 14365 27813 14399
rect 27813 14365 27847 14399
rect 27847 14365 27856 14399
rect 27804 14356 27856 14365
rect 20444 14220 20496 14272
rect 20536 14220 20588 14272
rect 22836 14220 22888 14272
rect 23296 14331 23348 14340
rect 23296 14297 23305 14331
rect 23305 14297 23339 14331
rect 23339 14297 23348 14331
rect 23296 14288 23348 14297
rect 24124 14288 24176 14340
rect 23848 14220 23900 14272
rect 24952 14263 25004 14272
rect 24952 14229 24961 14263
rect 24961 14229 24995 14263
rect 24995 14229 25004 14263
rect 24952 14220 25004 14229
rect 4874 14118 4926 14170
rect 4938 14118 4990 14170
rect 5002 14118 5054 14170
rect 5066 14118 5118 14170
rect 5130 14118 5182 14170
rect 2780 14059 2832 14068
rect 2780 14025 2789 14059
rect 2789 14025 2823 14059
rect 2823 14025 2832 14059
rect 2780 14016 2832 14025
rect 3240 13948 3292 14000
rect 1400 13923 1452 13932
rect 1400 13889 1409 13923
rect 1409 13889 1443 13923
rect 1443 13889 1452 13923
rect 1400 13880 1452 13889
rect 2688 13880 2740 13932
rect 3148 13923 3200 13932
rect 3148 13889 3157 13923
rect 3157 13889 3191 13923
rect 3191 13889 3200 13923
rect 3148 13880 3200 13889
rect 3608 14059 3660 14068
rect 3608 14025 3617 14059
rect 3617 14025 3651 14059
rect 3651 14025 3660 14059
rect 3608 14016 3660 14025
rect 3700 13923 3752 13932
rect 3700 13889 3709 13923
rect 3709 13889 3743 13923
rect 3743 13889 3752 13923
rect 3700 13880 3752 13889
rect 2320 13855 2372 13864
rect 2320 13821 2329 13855
rect 2329 13821 2363 13855
rect 2363 13821 2372 13855
rect 2320 13812 2372 13821
rect 2964 13855 3016 13864
rect 2964 13821 2973 13855
rect 2973 13821 3007 13855
rect 3007 13821 3016 13855
rect 2964 13812 3016 13821
rect 2228 13744 2280 13796
rect 4160 13923 4212 13932
rect 4160 13889 4169 13923
rect 4169 13889 4203 13923
rect 4203 13889 4212 13923
rect 4160 13880 4212 13889
rect 4252 13880 4304 13932
rect 4804 13880 4856 13932
rect 6736 13880 6788 13932
rect 5908 13855 5960 13864
rect 5908 13821 5917 13855
rect 5917 13821 5951 13855
rect 5951 13821 5960 13855
rect 5908 13812 5960 13821
rect 7012 13880 7064 13932
rect 7564 13923 7616 13932
rect 7564 13889 7573 13923
rect 7573 13889 7607 13923
rect 7607 13889 7616 13923
rect 7564 13880 7616 13889
rect 8300 13880 8352 13932
rect 9588 13923 9640 13932
rect 9588 13889 9597 13923
rect 9597 13889 9631 13923
rect 9631 13889 9640 13923
rect 9588 13880 9640 13889
rect 9680 13923 9732 13932
rect 9680 13889 9689 13923
rect 9689 13889 9723 13923
rect 9723 13889 9732 13923
rect 9680 13880 9732 13889
rect 11244 13880 11296 13932
rect 11888 13948 11940 14000
rect 13452 13991 13504 14000
rect 13452 13957 13461 13991
rect 13461 13957 13495 13991
rect 13495 13957 13504 13991
rect 13452 13948 13504 13957
rect 12900 13880 12952 13932
rect 13084 13880 13136 13932
rect 14096 13880 14148 13932
rect 16488 14016 16540 14068
rect 17132 14016 17184 14068
rect 14648 13991 14700 14000
rect 14648 13957 14657 13991
rect 14657 13957 14691 13991
rect 14691 13957 14700 13991
rect 14648 13948 14700 13957
rect 8668 13855 8720 13864
rect 8668 13821 8677 13855
rect 8677 13821 8711 13855
rect 8711 13821 8720 13855
rect 8668 13812 8720 13821
rect 16580 13948 16632 14000
rect 15936 13880 15988 13932
rect 18236 13948 18288 14000
rect 16856 13923 16908 13932
rect 16856 13889 16865 13923
rect 16865 13889 16899 13923
rect 16899 13889 16908 13923
rect 16856 13880 16908 13889
rect 18604 14016 18656 14068
rect 20536 14016 20588 14068
rect 20720 14016 20772 14068
rect 21548 14016 21600 14068
rect 18420 13948 18472 14000
rect 18880 13948 18932 14000
rect 17776 13812 17828 13864
rect 17960 13812 18012 13864
rect 6920 13744 6972 13796
rect 8576 13744 8628 13796
rect 13728 13744 13780 13796
rect 18788 13880 18840 13932
rect 18972 13923 19024 13932
rect 18972 13889 18981 13923
rect 18981 13889 19015 13923
rect 19015 13889 19024 13923
rect 18972 13880 19024 13889
rect 19156 13948 19208 14000
rect 19708 13880 19760 13932
rect 4620 13676 4672 13728
rect 9128 13719 9180 13728
rect 9128 13685 9137 13719
rect 9137 13685 9171 13719
rect 9171 13685 9180 13719
rect 9128 13676 9180 13685
rect 9220 13719 9272 13728
rect 9220 13685 9229 13719
rect 9229 13685 9263 13719
rect 9263 13685 9272 13719
rect 9220 13676 9272 13685
rect 12808 13676 12860 13728
rect 13820 13719 13872 13728
rect 13820 13685 13829 13719
rect 13829 13685 13863 13719
rect 13863 13685 13872 13719
rect 13820 13676 13872 13685
rect 14740 13676 14792 13728
rect 15384 13676 15436 13728
rect 18052 13676 18104 13728
rect 18880 13812 18932 13864
rect 20444 13812 20496 13864
rect 20536 13855 20588 13864
rect 20536 13821 20545 13855
rect 20545 13821 20579 13855
rect 20579 13821 20588 13855
rect 20536 13812 20588 13821
rect 20628 13855 20680 13864
rect 20628 13821 20637 13855
rect 20637 13821 20671 13855
rect 20671 13821 20680 13855
rect 20628 13812 20680 13821
rect 20904 13923 20956 13932
rect 20904 13889 20913 13923
rect 20913 13889 20947 13923
rect 20947 13889 20956 13923
rect 20904 13880 20956 13889
rect 21364 13948 21416 14000
rect 22376 13948 22428 14000
rect 21640 13923 21692 13932
rect 21640 13889 21649 13923
rect 21649 13889 21683 13923
rect 21683 13889 21692 13923
rect 21640 13880 21692 13889
rect 22284 13923 22336 13932
rect 22284 13889 22293 13923
rect 22293 13889 22327 13923
rect 22327 13889 22336 13923
rect 22284 13880 22336 13889
rect 22468 13923 22520 13932
rect 22468 13889 22477 13923
rect 22477 13889 22511 13923
rect 22511 13889 22520 13923
rect 22468 13880 22520 13889
rect 22560 13923 22612 13932
rect 22560 13889 22569 13923
rect 22569 13889 22603 13923
rect 22603 13889 22612 13923
rect 22560 13880 22612 13889
rect 23388 14016 23440 14068
rect 24584 14016 24636 14068
rect 23020 13923 23072 13932
rect 23020 13889 23029 13923
rect 23029 13889 23063 13923
rect 23063 13889 23072 13923
rect 23020 13880 23072 13889
rect 25228 13948 25280 14000
rect 23480 13880 23532 13932
rect 23572 13855 23624 13864
rect 23572 13821 23581 13855
rect 23581 13821 23615 13855
rect 23615 13821 23624 13855
rect 23572 13812 23624 13821
rect 23848 13855 23900 13864
rect 23848 13821 23857 13855
rect 23857 13821 23891 13855
rect 23891 13821 23900 13855
rect 23848 13812 23900 13821
rect 18604 13744 18656 13796
rect 18972 13676 19024 13728
rect 20260 13744 20312 13796
rect 22560 13744 22612 13796
rect 22928 13744 22980 13796
rect 19524 13676 19576 13728
rect 19616 13719 19668 13728
rect 19616 13685 19625 13719
rect 19625 13685 19659 13719
rect 19659 13685 19668 13719
rect 19616 13676 19668 13685
rect 19984 13676 20036 13728
rect 20352 13676 20404 13728
rect 23388 13676 23440 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 8760 13515 8812 13524
rect 8760 13481 8769 13515
rect 8769 13481 8803 13515
rect 8803 13481 8812 13515
rect 8760 13472 8812 13481
rect 10232 13515 10284 13524
rect 10232 13481 10241 13515
rect 10241 13481 10275 13515
rect 10275 13481 10284 13515
rect 10232 13472 10284 13481
rect 10416 13472 10468 13524
rect 13820 13472 13872 13524
rect 14832 13472 14884 13524
rect 15292 13472 15344 13524
rect 15568 13472 15620 13524
rect 15844 13472 15896 13524
rect 18972 13472 19024 13524
rect 19616 13472 19668 13524
rect 19708 13472 19760 13524
rect 20352 13472 20404 13524
rect 21364 13472 21416 13524
rect 2964 13379 3016 13388
rect 2964 13345 2973 13379
rect 2973 13345 3007 13379
rect 3007 13345 3016 13379
rect 2964 13336 3016 13345
rect 2688 13200 2740 13252
rect 3148 13268 3200 13320
rect 4712 13379 4764 13388
rect 4712 13345 4721 13379
rect 4721 13345 4755 13379
rect 4755 13345 4764 13379
rect 4712 13336 4764 13345
rect 8208 13404 8260 13456
rect 4620 13311 4672 13320
rect 4620 13277 4629 13311
rect 4629 13277 4663 13311
rect 4663 13277 4672 13311
rect 4620 13268 4672 13277
rect 6920 13311 6972 13320
rect 6920 13277 6929 13311
rect 6929 13277 6963 13311
rect 6963 13277 6972 13311
rect 6920 13268 6972 13277
rect 7012 13268 7064 13320
rect 8208 13311 8260 13320
rect 8208 13277 8217 13311
rect 8217 13277 8251 13311
rect 8251 13277 8260 13311
rect 8208 13268 8260 13277
rect 8668 13336 8720 13388
rect 9128 13379 9180 13388
rect 9128 13345 9137 13379
rect 9137 13345 9171 13379
rect 9171 13345 9180 13379
rect 9128 13336 9180 13345
rect 8484 13311 8536 13320
rect 8484 13277 8493 13311
rect 8493 13277 8527 13311
rect 8527 13277 8536 13311
rect 8484 13268 8536 13277
rect 7104 13243 7156 13252
rect 7104 13209 7113 13243
rect 7113 13209 7147 13243
rect 7147 13209 7156 13243
rect 7104 13200 7156 13209
rect 7564 13200 7616 13252
rect 9220 13311 9272 13320
rect 9220 13277 9229 13311
rect 9229 13277 9263 13311
rect 9263 13277 9272 13311
rect 9220 13268 9272 13277
rect 17040 13404 17092 13456
rect 12256 13336 12308 13388
rect 10232 13268 10284 13320
rect 12348 13268 12400 13320
rect 12716 13311 12768 13320
rect 12716 13277 12725 13311
rect 12725 13277 12759 13311
rect 12759 13277 12768 13311
rect 12716 13268 12768 13277
rect 12808 13311 12860 13320
rect 12808 13277 12817 13311
rect 12817 13277 12851 13311
rect 12851 13277 12860 13311
rect 12808 13268 12860 13277
rect 12992 13311 13044 13320
rect 12992 13277 13001 13311
rect 13001 13277 13035 13311
rect 13035 13277 13044 13311
rect 12992 13268 13044 13277
rect 9680 13200 9732 13252
rect 3792 13132 3844 13184
rect 5264 13175 5316 13184
rect 5264 13141 5273 13175
rect 5273 13141 5307 13175
rect 5307 13141 5316 13175
rect 5264 13132 5316 13141
rect 10048 13175 10100 13184
rect 10048 13141 10057 13175
rect 10057 13141 10091 13175
rect 10091 13141 10100 13175
rect 10048 13132 10100 13141
rect 11704 13243 11756 13252
rect 11704 13209 11713 13243
rect 11713 13209 11747 13243
rect 11747 13209 11756 13243
rect 11704 13200 11756 13209
rect 13912 13336 13964 13388
rect 14004 13336 14056 13388
rect 12164 13132 12216 13184
rect 12532 13132 12584 13184
rect 13544 13311 13596 13320
rect 13544 13277 13553 13311
rect 13553 13277 13587 13311
rect 13587 13277 13596 13311
rect 13544 13268 13596 13277
rect 14648 13311 14700 13320
rect 14648 13277 14657 13311
rect 14657 13277 14691 13311
rect 14691 13277 14700 13311
rect 14648 13268 14700 13277
rect 14924 13268 14976 13320
rect 15108 13311 15160 13320
rect 15108 13277 15117 13311
rect 15117 13277 15151 13311
rect 15151 13277 15160 13311
rect 15108 13268 15160 13277
rect 15292 13311 15344 13320
rect 15292 13277 15301 13311
rect 15301 13277 15335 13311
rect 15335 13277 15344 13311
rect 15292 13268 15344 13277
rect 15844 13379 15896 13388
rect 15844 13345 15853 13379
rect 15853 13345 15887 13379
rect 15887 13345 15896 13379
rect 15844 13336 15896 13345
rect 15936 13379 15988 13388
rect 15936 13345 15945 13379
rect 15945 13345 15979 13379
rect 15979 13345 15988 13379
rect 15936 13336 15988 13345
rect 15660 13311 15712 13320
rect 15660 13277 15669 13311
rect 15669 13277 15703 13311
rect 15703 13277 15712 13311
rect 15660 13268 15712 13277
rect 17960 13336 18012 13388
rect 18880 13336 18932 13388
rect 13360 13132 13412 13184
rect 14096 13132 14148 13184
rect 16396 13200 16448 13252
rect 18420 13311 18472 13320
rect 18420 13277 18429 13311
rect 18429 13277 18463 13311
rect 18463 13277 18472 13311
rect 19984 13336 20036 13388
rect 21180 13336 21232 13388
rect 21640 13472 21692 13524
rect 21732 13472 21784 13524
rect 22192 13472 22244 13524
rect 23296 13472 23348 13524
rect 23572 13472 23624 13524
rect 21824 13404 21876 13456
rect 18420 13268 18472 13277
rect 19616 13311 19668 13320
rect 19616 13277 19625 13311
rect 19625 13277 19659 13311
rect 19659 13277 19668 13311
rect 19616 13268 19668 13277
rect 19708 13311 19760 13320
rect 19708 13277 19717 13311
rect 19717 13277 19751 13311
rect 19751 13277 19760 13311
rect 19708 13268 19760 13277
rect 22744 13336 22796 13388
rect 18696 13200 18748 13252
rect 21364 13200 21416 13252
rect 21916 13200 21968 13252
rect 22100 13311 22152 13320
rect 22100 13277 22109 13311
rect 22109 13277 22143 13311
rect 22143 13277 22152 13311
rect 22100 13268 22152 13277
rect 22192 13311 22244 13320
rect 22192 13277 22201 13311
rect 22201 13277 22235 13311
rect 22235 13277 22244 13311
rect 22192 13268 22244 13277
rect 24952 13404 25004 13456
rect 22928 13379 22980 13388
rect 22928 13345 22937 13379
rect 22937 13345 22971 13379
rect 22971 13345 22980 13379
rect 22928 13336 22980 13345
rect 23204 13379 23256 13388
rect 23204 13345 23213 13379
rect 23213 13345 23247 13379
rect 23247 13345 23256 13379
rect 23204 13336 23256 13345
rect 24216 13268 24268 13320
rect 24584 13311 24636 13320
rect 24584 13277 24593 13311
rect 24593 13277 24627 13311
rect 24627 13277 24636 13311
rect 24584 13268 24636 13277
rect 22284 13200 22336 13252
rect 22560 13200 22612 13252
rect 24032 13200 24084 13252
rect 24768 13268 24820 13320
rect 16028 13132 16080 13184
rect 20260 13132 20312 13184
rect 21640 13132 21692 13184
rect 23756 13132 23808 13184
rect 4874 13030 4926 13082
rect 4938 13030 4990 13082
rect 5002 13030 5054 13082
rect 5066 13030 5118 13082
rect 5130 13030 5182 13082
rect 2228 12971 2280 12980
rect 2228 12937 2237 12971
rect 2237 12937 2271 12971
rect 2271 12937 2280 12971
rect 2228 12928 2280 12937
rect 5264 12928 5316 12980
rect 7104 12928 7156 12980
rect 8300 12928 8352 12980
rect 12716 12928 12768 12980
rect 16396 12928 16448 12980
rect 17776 12928 17828 12980
rect 18696 12971 18748 12980
rect 18696 12937 18705 12971
rect 18705 12937 18739 12971
rect 18739 12937 18748 12971
rect 18696 12928 18748 12937
rect 20168 12928 20220 12980
rect 22376 12928 22428 12980
rect 22744 12928 22796 12980
rect 2136 12792 2188 12844
rect 2412 12835 2464 12844
rect 2412 12801 2421 12835
rect 2421 12801 2455 12835
rect 2455 12801 2464 12835
rect 2412 12792 2464 12801
rect 4712 12792 4764 12844
rect 12992 12903 13044 12912
rect 12992 12869 13001 12903
rect 13001 12869 13035 12903
rect 13035 12869 13044 12903
rect 12992 12860 13044 12869
rect 14924 12860 14976 12912
rect 6184 12767 6236 12776
rect 6184 12733 6193 12767
rect 6193 12733 6227 12767
rect 6227 12733 6236 12767
rect 6184 12724 6236 12733
rect 7196 12835 7248 12844
rect 7196 12801 7205 12835
rect 7205 12801 7239 12835
rect 7239 12801 7248 12835
rect 7196 12792 7248 12801
rect 7472 12792 7524 12844
rect 8484 12792 8536 12844
rect 9588 12792 9640 12844
rect 15844 12860 15896 12912
rect 19800 12860 19852 12912
rect 20076 12903 20128 12912
rect 20076 12869 20085 12903
rect 20085 12869 20119 12903
rect 20119 12869 20128 12903
rect 20076 12860 20128 12869
rect 13544 12792 13596 12844
rect 14648 12792 14700 12844
rect 15384 12835 15436 12844
rect 15384 12801 15393 12835
rect 15393 12801 15427 12835
rect 15427 12801 15436 12835
rect 15384 12792 15436 12801
rect 15568 12835 15620 12844
rect 15568 12801 15577 12835
rect 15577 12801 15611 12835
rect 15611 12801 15620 12835
rect 15568 12792 15620 12801
rect 16120 12792 16172 12844
rect 18512 12792 18564 12844
rect 9680 12724 9732 12776
rect 10968 12724 11020 12776
rect 19616 12792 19668 12844
rect 19708 12835 19760 12844
rect 19708 12801 19717 12835
rect 19717 12801 19751 12835
rect 19751 12801 19760 12835
rect 19708 12792 19760 12801
rect 21640 12860 21692 12912
rect 22284 12860 22336 12912
rect 20352 12835 20404 12844
rect 20352 12801 20361 12835
rect 20361 12801 20395 12835
rect 20395 12801 20404 12835
rect 20352 12792 20404 12801
rect 20536 12792 20588 12844
rect 15844 12656 15896 12708
rect 20260 12724 20312 12776
rect 20812 12792 20864 12844
rect 20996 12835 21048 12844
rect 20996 12801 21005 12835
rect 21005 12801 21039 12835
rect 21039 12801 21048 12835
rect 20996 12792 21048 12801
rect 21180 12835 21232 12844
rect 21180 12801 21189 12835
rect 21189 12801 21223 12835
rect 21223 12801 21232 12835
rect 21180 12792 21232 12801
rect 22008 12835 22060 12844
rect 22008 12801 22017 12835
rect 22017 12801 22051 12835
rect 22051 12801 22060 12835
rect 22008 12792 22060 12801
rect 22836 12860 22888 12912
rect 22100 12724 22152 12776
rect 12808 12588 12860 12640
rect 13268 12588 13320 12640
rect 15292 12588 15344 12640
rect 15660 12588 15712 12640
rect 17040 12631 17092 12640
rect 17040 12597 17049 12631
rect 17049 12597 17083 12631
rect 17083 12597 17092 12631
rect 17040 12588 17092 12597
rect 19524 12588 19576 12640
rect 19892 12588 19944 12640
rect 20168 12588 20220 12640
rect 22192 12656 22244 12708
rect 23388 12835 23440 12844
rect 23388 12801 23397 12835
rect 23397 12801 23431 12835
rect 23431 12801 23440 12835
rect 23388 12792 23440 12801
rect 24032 12860 24084 12912
rect 24860 12928 24912 12980
rect 23572 12724 23624 12776
rect 20720 12631 20772 12640
rect 20720 12597 20729 12631
rect 20729 12597 20763 12631
rect 20763 12597 20772 12631
rect 20720 12588 20772 12597
rect 21088 12631 21140 12640
rect 21088 12597 21097 12631
rect 21097 12597 21131 12631
rect 21131 12597 21140 12631
rect 21088 12588 21140 12597
rect 23204 12631 23256 12640
rect 23204 12597 23213 12631
rect 23213 12597 23247 12631
rect 23247 12597 23256 12631
rect 23204 12588 23256 12597
rect 23296 12588 23348 12640
rect 24308 12588 24360 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 11152 12384 11204 12436
rect 15384 12384 15436 12436
rect 15844 12427 15896 12436
rect 1860 12316 1912 12368
rect 2688 12316 2740 12368
rect 13728 12316 13780 12368
rect 15844 12393 15853 12427
rect 15853 12393 15887 12427
rect 15887 12393 15896 12427
rect 15844 12384 15896 12393
rect 15936 12384 15988 12436
rect 2412 12291 2464 12300
rect 2412 12257 2421 12291
rect 2421 12257 2455 12291
rect 2455 12257 2464 12291
rect 2412 12248 2464 12257
rect 6184 12248 6236 12300
rect 7472 12291 7524 12300
rect 7472 12257 7481 12291
rect 7481 12257 7515 12291
rect 7515 12257 7524 12291
rect 7472 12248 7524 12257
rect 12900 12248 12952 12300
rect 14096 12248 14148 12300
rect 15844 12248 15896 12300
rect 19432 12384 19484 12436
rect 16580 12316 16632 12368
rect 17684 12316 17736 12368
rect 18696 12316 18748 12368
rect 2044 12180 2096 12232
rect 2136 12180 2188 12232
rect 8484 12180 8536 12232
rect 12532 12223 12584 12232
rect 12532 12189 12541 12223
rect 12541 12189 12575 12223
rect 12575 12189 12584 12223
rect 12532 12180 12584 12189
rect 12624 12223 12676 12232
rect 12624 12189 12633 12223
rect 12633 12189 12667 12223
rect 12667 12189 12676 12223
rect 12624 12180 12676 12189
rect 13176 12180 13228 12232
rect 12716 12112 12768 12164
rect 16856 12248 16908 12300
rect 20720 12248 20772 12300
rect 15384 12155 15436 12164
rect 15384 12121 15393 12155
rect 15393 12121 15427 12155
rect 15427 12121 15436 12155
rect 15384 12112 15436 12121
rect 15568 12155 15620 12164
rect 15568 12121 15593 12155
rect 15593 12121 15620 12155
rect 15568 12112 15620 12121
rect 15844 12155 15896 12164
rect 15844 12121 15853 12155
rect 15853 12121 15887 12155
rect 15887 12121 15896 12155
rect 15844 12112 15896 12121
rect 16488 12180 16540 12232
rect 19340 12180 19392 12232
rect 16580 12112 16632 12164
rect 16948 12112 17000 12164
rect 2872 12087 2924 12096
rect 2872 12053 2881 12087
rect 2881 12053 2915 12087
rect 2915 12053 2924 12087
rect 2872 12044 2924 12053
rect 7012 12044 7064 12096
rect 15936 12044 15988 12096
rect 18420 12044 18472 12096
rect 19800 12180 19852 12232
rect 21088 12180 21140 12232
rect 19524 12112 19576 12164
rect 21272 12112 21324 12164
rect 20536 12044 20588 12096
rect 23480 12044 23532 12096
rect 24676 12044 24728 12096
rect 4874 11942 4926 11994
rect 4938 11942 4990 11994
rect 5002 11942 5054 11994
rect 5066 11942 5118 11994
rect 5130 11942 5182 11994
rect 848 11704 900 11756
rect 4528 11840 4580 11892
rect 12440 11840 12492 11892
rect 12624 11840 12676 11892
rect 12992 11840 13044 11892
rect 13176 11883 13228 11892
rect 13176 11849 13185 11883
rect 13185 11849 13219 11883
rect 13219 11849 13228 11883
rect 13176 11840 13228 11849
rect 13360 11840 13412 11892
rect 4712 11815 4764 11824
rect 4712 11781 4721 11815
rect 4721 11781 4755 11815
rect 4755 11781 4764 11815
rect 4712 11772 4764 11781
rect 4804 11772 4856 11824
rect 1952 11636 2004 11688
rect 3792 11679 3844 11688
rect 3792 11645 3801 11679
rect 3801 11645 3835 11679
rect 3835 11645 3844 11679
rect 7656 11772 7708 11824
rect 4528 11747 4580 11756
rect 4528 11713 4537 11747
rect 4537 11713 4571 11747
rect 4571 11713 4580 11747
rect 4528 11704 4580 11713
rect 4896 11747 4948 11756
rect 3792 11636 3844 11645
rect 4896 11713 4905 11747
rect 4905 11713 4939 11747
rect 4939 11713 4948 11747
rect 4896 11704 4948 11713
rect 5356 11747 5408 11756
rect 5356 11713 5365 11747
rect 5365 11713 5399 11747
rect 5399 11713 5408 11747
rect 5356 11704 5408 11713
rect 5540 11636 5592 11688
rect 8760 11747 8812 11756
rect 8760 11713 8769 11747
rect 8769 11713 8803 11747
rect 8803 11713 8812 11747
rect 8760 11704 8812 11713
rect 10968 11815 11020 11824
rect 10968 11781 10977 11815
rect 10977 11781 11011 11815
rect 11011 11781 11020 11815
rect 10968 11772 11020 11781
rect 11060 11772 11112 11824
rect 9220 11636 9272 11688
rect 9864 11747 9916 11756
rect 9864 11713 9873 11747
rect 9873 11713 9907 11747
rect 9907 11713 9916 11747
rect 9864 11704 9916 11713
rect 10232 11704 10284 11756
rect 12256 11704 12308 11756
rect 9772 11636 9824 11688
rect 8760 11568 8812 11620
rect 11336 11611 11388 11620
rect 11336 11577 11345 11611
rect 11345 11577 11379 11611
rect 11379 11577 11388 11611
rect 11336 11568 11388 11577
rect 12624 11636 12676 11688
rect 13084 11747 13136 11756
rect 13084 11713 13093 11747
rect 13093 11713 13127 11747
rect 13127 11713 13136 11747
rect 13084 11704 13136 11713
rect 13176 11704 13228 11756
rect 13912 11772 13964 11824
rect 14648 11840 14700 11892
rect 13820 11747 13872 11756
rect 13820 11713 13829 11747
rect 13829 11713 13863 11747
rect 13863 11713 13872 11747
rect 13820 11704 13872 11713
rect 13728 11636 13780 11688
rect 15476 11840 15528 11892
rect 15568 11883 15620 11892
rect 15568 11849 15577 11883
rect 15577 11849 15611 11883
rect 15611 11849 15620 11883
rect 15568 11840 15620 11849
rect 19340 11840 19392 11892
rect 19984 11883 20036 11892
rect 19984 11849 19993 11883
rect 19993 11849 20027 11883
rect 20027 11849 20036 11883
rect 19984 11840 20036 11849
rect 20168 11840 20220 11892
rect 15568 11704 15620 11756
rect 15936 11747 15988 11756
rect 15936 11713 15945 11747
rect 15945 11713 15979 11747
rect 15979 11713 15988 11747
rect 15936 11704 15988 11713
rect 15476 11679 15528 11688
rect 15476 11645 15485 11679
rect 15485 11645 15519 11679
rect 15519 11645 15528 11679
rect 15476 11636 15528 11645
rect 22652 11772 22704 11824
rect 23572 11840 23624 11892
rect 25136 11840 25188 11892
rect 24400 11772 24452 11824
rect 16120 11747 16172 11756
rect 16120 11713 16129 11747
rect 16129 11713 16163 11747
rect 16163 11713 16172 11747
rect 16120 11704 16172 11713
rect 16304 11747 16356 11756
rect 16304 11713 16313 11747
rect 16313 11713 16347 11747
rect 16347 11713 16356 11747
rect 16304 11704 16356 11713
rect 9588 11500 9640 11552
rect 11152 11543 11204 11552
rect 11152 11509 11161 11543
rect 11161 11509 11195 11543
rect 11195 11509 11204 11543
rect 11152 11500 11204 11509
rect 13176 11500 13228 11552
rect 13452 11500 13504 11552
rect 13544 11500 13596 11552
rect 13820 11500 13872 11552
rect 14464 11500 14516 11552
rect 15200 11500 15252 11552
rect 16028 11500 16080 11552
rect 16488 11704 16540 11756
rect 17224 11704 17276 11756
rect 18420 11747 18472 11756
rect 18420 11713 18429 11747
rect 18429 11713 18463 11747
rect 18463 11713 18472 11747
rect 18420 11704 18472 11713
rect 17040 11568 17092 11620
rect 16764 11500 16816 11552
rect 16948 11500 17000 11552
rect 18604 11500 18656 11552
rect 18788 11543 18840 11552
rect 18788 11509 18797 11543
rect 18797 11509 18831 11543
rect 18831 11509 18840 11543
rect 18788 11500 18840 11509
rect 19616 11679 19668 11688
rect 19616 11645 19625 11679
rect 19625 11645 19659 11679
rect 19659 11645 19668 11679
rect 19616 11636 19668 11645
rect 21088 11704 21140 11756
rect 23848 11747 23900 11756
rect 23848 11713 23857 11747
rect 23857 11713 23891 11747
rect 23891 11713 23900 11747
rect 23848 11704 23900 11713
rect 24124 11704 24176 11756
rect 19984 11500 20036 11552
rect 20812 11636 20864 11688
rect 24308 11747 24360 11756
rect 24308 11713 24317 11747
rect 24317 11713 24351 11747
rect 24351 11713 24360 11747
rect 24308 11704 24360 11713
rect 24860 11704 24912 11756
rect 25688 11747 25740 11756
rect 25688 11713 25697 11747
rect 25697 11713 25731 11747
rect 25731 11713 25740 11747
rect 25688 11704 25740 11713
rect 26608 11704 26660 11756
rect 24492 11636 24544 11688
rect 20720 11500 20772 11552
rect 24032 11500 24084 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 4620 11296 4672 11348
rect 11060 11296 11112 11348
rect 12164 11339 12216 11348
rect 12164 11305 12173 11339
rect 12173 11305 12207 11339
rect 12207 11305 12216 11339
rect 12164 11296 12216 11305
rect 12532 11296 12584 11348
rect 13176 11339 13228 11348
rect 13176 11305 13185 11339
rect 13185 11305 13219 11339
rect 13219 11305 13228 11339
rect 13176 11296 13228 11305
rect 13636 11296 13688 11348
rect 15844 11296 15896 11348
rect 4804 11160 4856 11212
rect 4896 11203 4948 11212
rect 4896 11169 4905 11203
rect 4905 11169 4939 11203
rect 4939 11169 4948 11203
rect 4896 11160 4948 11169
rect 2872 11092 2924 11144
rect 3148 11135 3200 11144
rect 3148 11101 3157 11135
rect 3157 11101 3191 11135
rect 3191 11101 3200 11135
rect 3148 11092 3200 11101
rect 1952 11024 2004 11076
rect 4160 11135 4212 11144
rect 4160 11101 4169 11135
rect 4169 11101 4203 11135
rect 4203 11101 4212 11135
rect 4160 11092 4212 11101
rect 7196 11271 7248 11280
rect 7196 11237 7205 11271
rect 7205 11237 7239 11271
rect 7239 11237 7248 11271
rect 7196 11228 7248 11237
rect 11428 11228 11480 11280
rect 5356 11160 5408 11212
rect 5540 11092 5592 11144
rect 7564 11203 7616 11212
rect 7564 11169 7573 11203
rect 7573 11169 7607 11203
rect 7607 11169 7616 11203
rect 7564 11160 7616 11169
rect 11612 11160 11664 11212
rect 8576 11092 8628 11144
rect 9588 11092 9640 11144
rect 9772 11092 9824 11144
rect 9956 11092 10008 11144
rect 10600 11135 10652 11144
rect 10600 11101 10609 11135
rect 10609 11101 10643 11135
rect 10643 11101 10652 11135
rect 10600 11092 10652 11101
rect 11520 11092 11572 11144
rect 11888 11160 11940 11212
rect 12900 11228 12952 11280
rect 15476 11228 15528 11280
rect 15936 11228 15988 11280
rect 11980 11135 12032 11144
rect 11980 11101 11989 11135
rect 11989 11101 12023 11135
rect 12023 11101 12032 11135
rect 11980 11092 12032 11101
rect 12348 11092 12400 11144
rect 12716 11092 12768 11144
rect 13084 11203 13136 11212
rect 13084 11169 13093 11203
rect 13093 11169 13127 11203
rect 13127 11169 13136 11203
rect 13084 11160 13136 11169
rect 13636 11160 13688 11212
rect 15200 11160 15252 11212
rect 16396 11296 16448 11348
rect 17224 11296 17276 11348
rect 18696 11296 18748 11348
rect 19800 11339 19852 11348
rect 19800 11305 19809 11339
rect 19809 11305 19843 11339
rect 19843 11305 19852 11339
rect 19800 11296 19852 11305
rect 19984 11296 20036 11348
rect 21180 11296 21232 11348
rect 21364 11296 21416 11348
rect 21548 11296 21600 11348
rect 17684 11228 17736 11280
rect 20168 11228 20220 11280
rect 13268 11135 13320 11144
rect 13268 11101 13277 11135
rect 13277 11101 13311 11135
rect 13311 11101 13320 11135
rect 13268 11092 13320 11101
rect 13544 11135 13596 11144
rect 13544 11101 13553 11135
rect 13553 11101 13587 11135
rect 13587 11101 13596 11135
rect 13544 11092 13596 11101
rect 13728 11135 13780 11144
rect 13728 11101 13737 11135
rect 13737 11101 13771 11135
rect 13771 11101 13780 11135
rect 13728 11092 13780 11101
rect 15384 11135 15436 11144
rect 15384 11101 15393 11135
rect 15393 11101 15427 11135
rect 15427 11101 15436 11135
rect 15384 11092 15436 11101
rect 5816 11024 5868 11076
rect 4712 10956 4764 11008
rect 6460 10956 6512 11008
rect 6736 10956 6788 11008
rect 8668 10956 8720 11008
rect 10692 11067 10744 11076
rect 10692 11033 10701 11067
rect 10701 11033 10735 11067
rect 10735 11033 10744 11067
rect 10692 11024 10744 11033
rect 10876 11067 10928 11076
rect 10876 11033 10885 11067
rect 10885 11033 10919 11067
rect 10919 11033 10928 11067
rect 10876 11024 10928 11033
rect 14004 11024 14056 11076
rect 15660 11135 15712 11144
rect 15660 11101 15669 11135
rect 15669 11101 15703 11135
rect 15703 11101 15712 11135
rect 15660 11092 15712 11101
rect 15752 11092 15804 11144
rect 16948 11160 17000 11212
rect 16028 11135 16080 11144
rect 16028 11101 16037 11135
rect 16037 11101 16071 11135
rect 16071 11101 16080 11135
rect 16028 11092 16080 11101
rect 16212 11092 16264 11144
rect 18328 11135 18380 11144
rect 18328 11101 18337 11135
rect 18337 11101 18371 11135
rect 18371 11101 18380 11135
rect 18328 11092 18380 11101
rect 19340 11135 19392 11144
rect 19340 11101 19349 11135
rect 19349 11101 19383 11135
rect 19383 11101 19392 11135
rect 19340 11092 19392 11101
rect 19432 11135 19484 11144
rect 19432 11101 19441 11135
rect 19441 11101 19475 11135
rect 19475 11101 19484 11135
rect 19432 11092 19484 11101
rect 16488 11024 16540 11076
rect 18512 11067 18564 11076
rect 18512 11033 18521 11067
rect 18521 11033 18555 11067
rect 18555 11033 18564 11067
rect 18512 11024 18564 11033
rect 18972 11024 19024 11076
rect 19800 11092 19852 11144
rect 20444 11092 20496 11144
rect 21548 11203 21600 11212
rect 21548 11169 21557 11203
rect 21557 11169 21591 11203
rect 21591 11169 21600 11203
rect 21548 11160 21600 11169
rect 21272 11135 21324 11144
rect 21272 11101 21281 11135
rect 21281 11101 21315 11135
rect 21315 11101 21324 11135
rect 21272 11092 21324 11101
rect 21364 11135 21416 11144
rect 21364 11101 21373 11135
rect 21373 11101 21407 11135
rect 21407 11101 21416 11135
rect 21364 11092 21416 11101
rect 20812 11024 20864 11076
rect 23204 11135 23256 11144
rect 23204 11101 23213 11135
rect 23213 11101 23247 11135
rect 23247 11101 23256 11135
rect 23204 11092 23256 11101
rect 23664 11092 23716 11144
rect 24492 11296 24544 11348
rect 24860 11296 24912 11348
rect 23940 11228 23992 11280
rect 24676 11160 24728 11212
rect 23940 11135 23992 11144
rect 23940 11101 23949 11135
rect 23949 11101 23983 11135
rect 23983 11101 23992 11135
rect 23940 11092 23992 11101
rect 11980 10956 12032 11008
rect 12348 10956 12400 11008
rect 12624 10956 12676 11008
rect 12992 10956 13044 11008
rect 16120 10956 16172 11008
rect 16580 10956 16632 11008
rect 17592 10956 17644 11008
rect 20720 10956 20772 11008
rect 24216 11024 24268 11076
rect 24768 11024 24820 11076
rect 25136 11024 25188 11076
rect 24032 10956 24084 11008
rect 4874 10854 4926 10906
rect 4938 10854 4990 10906
rect 5002 10854 5054 10906
rect 5066 10854 5118 10906
rect 5130 10854 5182 10906
rect 3148 10752 3200 10804
rect 5816 10795 5868 10804
rect 5816 10761 5825 10795
rect 5825 10761 5859 10795
rect 5859 10761 5868 10795
rect 5816 10752 5868 10761
rect 8668 10795 8720 10804
rect 8668 10761 8677 10795
rect 8677 10761 8711 10795
rect 8711 10761 8720 10795
rect 8668 10752 8720 10761
rect 9864 10752 9916 10804
rect 1860 10659 1912 10668
rect 1860 10625 1869 10659
rect 1869 10625 1903 10659
rect 1903 10625 1912 10659
rect 1860 10616 1912 10625
rect 1952 10591 2004 10600
rect 1952 10557 1961 10591
rect 1961 10557 1995 10591
rect 1995 10557 2004 10591
rect 1952 10548 2004 10557
rect 2872 10548 2924 10600
rect 2688 10480 2740 10532
rect 3424 10616 3476 10668
rect 6460 10684 6512 10736
rect 8484 10684 8536 10736
rect 6368 10616 6420 10668
rect 8576 10659 8628 10668
rect 8576 10625 8585 10659
rect 8585 10625 8619 10659
rect 8619 10625 8628 10659
rect 8576 10616 8628 10625
rect 9772 10684 9824 10736
rect 9220 10659 9272 10668
rect 9220 10625 9229 10659
rect 9229 10625 9263 10659
rect 9263 10625 9272 10659
rect 9220 10616 9272 10625
rect 9864 10659 9916 10668
rect 9864 10625 9873 10659
rect 9873 10625 9907 10659
rect 9907 10625 9916 10659
rect 9864 10616 9916 10625
rect 6460 10591 6512 10600
rect 6460 10557 6469 10591
rect 6469 10557 6503 10591
rect 6503 10557 6512 10591
rect 6460 10548 6512 10557
rect 7564 10548 7616 10600
rect 8392 10548 8444 10600
rect 8852 10480 8904 10532
rect 10416 10616 10468 10668
rect 11520 10659 11572 10668
rect 11520 10625 11529 10659
rect 11529 10625 11563 10659
rect 11563 10625 11572 10659
rect 11520 10616 11572 10625
rect 11428 10548 11480 10600
rect 11796 10659 11848 10668
rect 11796 10625 11805 10659
rect 11805 10625 11839 10659
rect 11839 10625 11848 10659
rect 11796 10616 11848 10625
rect 11888 10659 11940 10668
rect 11888 10625 11897 10659
rect 11897 10625 11931 10659
rect 11931 10625 11940 10659
rect 11888 10616 11940 10625
rect 11980 10616 12032 10668
rect 12164 10659 12216 10668
rect 12164 10625 12173 10659
rect 12173 10625 12207 10659
rect 12207 10625 12216 10659
rect 12164 10616 12216 10625
rect 12624 10659 12676 10668
rect 12624 10625 12633 10659
rect 12633 10625 12667 10659
rect 12667 10625 12676 10659
rect 12624 10616 12676 10625
rect 12808 10659 12860 10668
rect 12808 10625 12817 10659
rect 12817 10625 12851 10659
rect 12851 10625 12860 10659
rect 12808 10616 12860 10625
rect 12992 10659 13044 10668
rect 12992 10625 13001 10659
rect 13001 10625 13035 10659
rect 13035 10625 13044 10659
rect 12992 10616 13044 10625
rect 15476 10795 15528 10804
rect 15476 10761 15485 10795
rect 15485 10761 15519 10795
rect 15519 10761 15528 10795
rect 15476 10752 15528 10761
rect 16304 10752 16356 10804
rect 18144 10795 18196 10804
rect 18144 10761 18153 10795
rect 18153 10761 18187 10795
rect 18187 10761 18196 10795
rect 18144 10752 18196 10761
rect 18420 10752 18472 10804
rect 18788 10752 18840 10804
rect 15936 10684 15988 10736
rect 14004 10659 14056 10668
rect 14004 10625 14013 10659
rect 14013 10625 14047 10659
rect 14047 10625 14056 10659
rect 14004 10616 14056 10625
rect 13268 10548 13320 10600
rect 14464 10659 14516 10668
rect 14464 10625 14473 10659
rect 14473 10625 14507 10659
rect 14507 10625 14516 10659
rect 14464 10616 14516 10625
rect 14740 10616 14792 10668
rect 16120 10616 16172 10668
rect 10692 10480 10744 10532
rect 14096 10480 14148 10532
rect 4068 10412 4120 10464
rect 5356 10412 5408 10464
rect 10416 10412 10468 10464
rect 12624 10412 12676 10464
rect 13452 10412 13504 10464
rect 15476 10548 15528 10600
rect 16304 10616 16356 10668
rect 16672 10659 16724 10668
rect 16672 10625 16681 10659
rect 16681 10625 16715 10659
rect 16715 10625 16724 10659
rect 16672 10616 16724 10625
rect 18512 10684 18564 10736
rect 23848 10752 23900 10804
rect 24492 10795 24544 10804
rect 24492 10761 24517 10795
rect 24517 10761 24544 10795
rect 24492 10752 24544 10761
rect 17224 10659 17276 10668
rect 17224 10625 17233 10659
rect 17233 10625 17267 10659
rect 17267 10625 17276 10659
rect 17224 10616 17276 10625
rect 17500 10659 17552 10668
rect 17500 10625 17509 10659
rect 17509 10625 17543 10659
rect 17543 10625 17552 10659
rect 17500 10616 17552 10625
rect 17592 10659 17644 10668
rect 17592 10625 17602 10659
rect 17602 10625 17636 10659
rect 17636 10625 17644 10659
rect 17592 10616 17644 10625
rect 17776 10659 17828 10668
rect 17776 10625 17785 10659
rect 17785 10625 17819 10659
rect 17819 10625 17828 10659
rect 17776 10616 17828 10625
rect 17868 10659 17920 10668
rect 17868 10625 17877 10659
rect 17877 10625 17911 10659
rect 17911 10625 17920 10659
rect 17868 10616 17920 10625
rect 18144 10616 18196 10668
rect 19892 10616 19944 10668
rect 20720 10616 20772 10668
rect 21180 10659 21232 10668
rect 21180 10625 21189 10659
rect 21189 10625 21223 10659
rect 21223 10625 21232 10659
rect 21180 10616 21232 10625
rect 21732 10684 21784 10736
rect 23756 10727 23808 10736
rect 23756 10693 23765 10727
rect 23765 10693 23799 10727
rect 23799 10693 23808 10727
rect 23756 10684 23808 10693
rect 24124 10684 24176 10736
rect 24400 10684 24452 10736
rect 21548 10659 21600 10668
rect 21548 10625 21557 10659
rect 21557 10625 21591 10659
rect 21591 10625 21600 10659
rect 21548 10616 21600 10625
rect 24032 10659 24084 10668
rect 24032 10625 24041 10659
rect 24041 10625 24075 10659
rect 24075 10625 24084 10659
rect 24032 10616 24084 10625
rect 14464 10412 14516 10464
rect 16028 10412 16080 10464
rect 16396 10412 16448 10464
rect 21824 10548 21876 10600
rect 21916 10548 21968 10600
rect 18604 10480 18656 10532
rect 20904 10480 20956 10532
rect 21732 10480 21784 10532
rect 23664 10480 23716 10532
rect 24584 10616 24636 10668
rect 24768 10480 24820 10532
rect 20260 10455 20312 10464
rect 20260 10421 20269 10455
rect 20269 10421 20303 10455
rect 20303 10421 20312 10455
rect 20260 10412 20312 10421
rect 23204 10412 23256 10464
rect 23848 10455 23900 10464
rect 23848 10421 23857 10455
rect 23857 10421 23891 10455
rect 23891 10421 23900 10455
rect 23848 10412 23900 10421
rect 24400 10412 24452 10464
rect 24952 10412 25004 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 8392 10208 8444 10260
rect 4620 10140 4672 10192
rect 2688 10115 2740 10124
rect 2688 10081 2697 10115
rect 2697 10081 2731 10115
rect 2731 10081 2740 10115
rect 2688 10072 2740 10081
rect 4068 10115 4120 10124
rect 4068 10081 4077 10115
rect 4077 10081 4111 10115
rect 4111 10081 4120 10115
rect 4068 10072 4120 10081
rect 3424 10004 3476 10056
rect 5356 10072 5408 10124
rect 5448 10072 5500 10124
rect 8300 10140 8352 10192
rect 8668 10208 8720 10260
rect 11888 10208 11940 10260
rect 12992 10251 13044 10260
rect 12992 10217 13001 10251
rect 13001 10217 13035 10251
rect 13035 10217 13044 10251
rect 12992 10208 13044 10217
rect 13084 10208 13136 10260
rect 13268 10208 13320 10260
rect 14740 10251 14792 10260
rect 14740 10217 14749 10251
rect 14749 10217 14783 10251
rect 14783 10217 14792 10251
rect 14740 10208 14792 10217
rect 16396 10251 16448 10260
rect 16396 10217 16405 10251
rect 16405 10217 16439 10251
rect 16439 10217 16448 10251
rect 16396 10208 16448 10217
rect 16672 10208 16724 10260
rect 22192 10208 22244 10260
rect 24492 10251 24544 10260
rect 24492 10217 24501 10251
rect 24501 10217 24535 10251
rect 24535 10217 24544 10251
rect 24492 10208 24544 10217
rect 24768 10208 24820 10260
rect 4712 10004 4764 10056
rect 5540 10004 5592 10056
rect 6736 10004 6788 10056
rect 8852 10072 8904 10124
rect 4804 9868 4856 9920
rect 8392 10047 8444 10056
rect 8392 10013 8401 10047
rect 8401 10013 8435 10047
rect 8435 10013 8444 10047
rect 8392 10004 8444 10013
rect 9036 10004 9088 10056
rect 9496 10047 9548 10056
rect 9496 10013 9505 10047
rect 9505 10013 9539 10047
rect 9539 10013 9548 10047
rect 9496 10004 9548 10013
rect 9680 10004 9732 10056
rect 11612 10047 11664 10056
rect 11612 10013 11621 10047
rect 11621 10013 11655 10047
rect 11655 10013 11664 10047
rect 11612 10004 11664 10013
rect 13544 10140 13596 10192
rect 14096 10140 14148 10192
rect 12164 10072 12216 10124
rect 14004 10072 14056 10124
rect 8300 9936 8352 9988
rect 9588 9979 9640 9988
rect 9588 9945 9597 9979
rect 9597 9945 9631 9979
rect 9631 9945 9640 9979
rect 9588 9936 9640 9945
rect 8760 9868 8812 9920
rect 11152 9936 11204 9988
rect 11520 9936 11572 9988
rect 12072 10004 12124 10056
rect 12624 10004 12676 10056
rect 12716 10047 12768 10056
rect 12716 10013 12725 10047
rect 12725 10013 12759 10047
rect 12759 10013 12768 10047
rect 12716 10004 12768 10013
rect 12900 10004 12952 10056
rect 13452 10047 13504 10056
rect 13452 10013 13461 10047
rect 13461 10013 13495 10047
rect 13495 10013 13504 10047
rect 13452 10004 13504 10013
rect 13544 10047 13596 10056
rect 13544 10013 13553 10047
rect 13553 10013 13587 10047
rect 13587 10013 13596 10047
rect 13544 10004 13596 10013
rect 14372 10047 14424 10056
rect 14372 10013 14381 10047
rect 14381 10013 14415 10047
rect 14415 10013 14424 10047
rect 14372 10004 14424 10013
rect 16764 10140 16816 10192
rect 17776 10140 17828 10192
rect 18328 10140 18380 10192
rect 19616 10140 19668 10192
rect 17224 10072 17276 10124
rect 17408 10072 17460 10124
rect 18144 10072 18196 10124
rect 19432 10072 19484 10124
rect 16580 10004 16632 10056
rect 16948 10004 17000 10056
rect 11428 9868 11480 9920
rect 14096 9979 14148 9988
rect 14096 9945 14105 9979
rect 14105 9945 14139 9979
rect 14139 9945 14148 9979
rect 14096 9936 14148 9945
rect 15476 9936 15528 9988
rect 18328 10047 18380 10056
rect 18328 10013 18337 10047
rect 18337 10013 18371 10047
rect 18371 10013 18380 10047
rect 18328 10004 18380 10013
rect 18788 10047 18840 10056
rect 18788 10013 18797 10047
rect 18797 10013 18831 10047
rect 18831 10013 18840 10047
rect 18788 10004 18840 10013
rect 20260 10072 20312 10124
rect 12164 9868 12216 9920
rect 12624 9911 12676 9920
rect 12624 9877 12633 9911
rect 12633 9877 12667 9911
rect 12667 9877 12676 9911
rect 12624 9868 12676 9877
rect 12716 9868 12768 9920
rect 13912 9868 13964 9920
rect 16304 9868 16356 9920
rect 17408 9936 17460 9988
rect 19064 9936 19116 9988
rect 19616 9979 19668 9988
rect 19616 9945 19625 9979
rect 19625 9945 19659 9979
rect 19659 9945 19668 9979
rect 19616 9936 19668 9945
rect 20168 10047 20220 10056
rect 20168 10013 20177 10047
rect 20177 10013 20211 10047
rect 20211 10013 20220 10047
rect 20168 10004 20220 10013
rect 20352 10004 20404 10056
rect 20536 10047 20588 10056
rect 20536 10013 20545 10047
rect 20545 10013 20579 10047
rect 20579 10013 20588 10047
rect 20536 10004 20588 10013
rect 24032 10004 24084 10056
rect 24952 10140 25004 10192
rect 24676 10072 24728 10124
rect 24584 10047 24636 10056
rect 24584 10013 24593 10047
rect 24593 10013 24627 10047
rect 24627 10013 24636 10047
rect 24584 10004 24636 10013
rect 19800 9868 19852 9920
rect 20812 9936 20864 9988
rect 21456 9936 21508 9988
rect 23572 9936 23624 9988
rect 20720 9868 20772 9920
rect 25044 9936 25096 9988
rect 25136 9868 25188 9920
rect 4874 9766 4926 9818
rect 4938 9766 4990 9818
rect 5002 9766 5054 9818
rect 5066 9766 5118 9818
rect 5130 9766 5182 9818
rect 9588 9664 9640 9716
rect 11152 9664 11204 9716
rect 8852 9596 8904 9648
rect 9496 9596 9548 9648
rect 12164 9571 12216 9580
rect 12164 9537 12173 9571
rect 12173 9537 12207 9571
rect 12207 9537 12216 9571
rect 12164 9528 12216 9537
rect 12256 9571 12308 9580
rect 12256 9537 12265 9571
rect 12265 9537 12299 9571
rect 12299 9537 12308 9571
rect 12256 9528 12308 9537
rect 12624 9528 12676 9580
rect 12992 9528 13044 9580
rect 13728 9596 13780 9648
rect 13452 9571 13504 9580
rect 13452 9537 13461 9571
rect 13461 9537 13495 9571
rect 13495 9537 13504 9571
rect 13452 9528 13504 9537
rect 13544 9528 13596 9580
rect 12716 9392 12768 9444
rect 12900 9392 12952 9444
rect 13636 9392 13688 9444
rect 18788 9664 18840 9716
rect 21456 9664 21508 9716
rect 19064 9596 19116 9648
rect 20812 9596 20864 9648
rect 18144 9571 18196 9580
rect 18144 9537 18153 9571
rect 18153 9537 18187 9571
rect 18187 9537 18196 9571
rect 18144 9528 18196 9537
rect 18236 9503 18288 9512
rect 18236 9469 18245 9503
rect 18245 9469 18279 9503
rect 18279 9469 18288 9503
rect 20168 9528 20220 9580
rect 21824 9707 21876 9716
rect 21824 9673 21833 9707
rect 21833 9673 21867 9707
rect 21867 9673 21876 9707
rect 21824 9664 21876 9673
rect 25044 9664 25096 9716
rect 22284 9596 22336 9648
rect 22192 9571 22244 9580
rect 22192 9537 22201 9571
rect 22201 9537 22235 9571
rect 22235 9537 22244 9571
rect 22192 9528 22244 9537
rect 22560 9571 22612 9580
rect 22560 9537 22569 9571
rect 22569 9537 22603 9571
rect 22603 9537 22612 9571
rect 22560 9528 22612 9537
rect 24032 9571 24084 9580
rect 24032 9537 24041 9571
rect 24041 9537 24075 9571
rect 24075 9537 24084 9571
rect 24032 9528 24084 9537
rect 24584 9528 24636 9580
rect 18236 9460 18288 9469
rect 18880 9460 18932 9512
rect 22376 9503 22428 9512
rect 22376 9469 22385 9503
rect 22385 9469 22419 9503
rect 22419 9469 22428 9503
rect 22376 9460 22428 9469
rect 18972 9435 19024 9444
rect 18972 9401 18981 9435
rect 18981 9401 19015 9435
rect 19015 9401 19024 9435
rect 18972 9392 19024 9401
rect 22008 9392 22060 9444
rect 8944 9367 8996 9376
rect 8944 9333 8953 9367
rect 8953 9333 8987 9367
rect 8987 9333 8996 9367
rect 8944 9324 8996 9333
rect 12256 9324 12308 9376
rect 12348 9324 12400 9376
rect 13268 9324 13320 9376
rect 17868 9324 17920 9376
rect 19616 9324 19668 9376
rect 19984 9324 20036 9376
rect 20720 9324 20772 9376
rect 21088 9367 21140 9376
rect 21088 9333 21097 9367
rect 21097 9333 21131 9367
rect 21131 9333 21140 9367
rect 21088 9324 21140 9333
rect 23664 9324 23716 9376
rect 24860 9324 24912 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 6276 9163 6328 9172
rect 6276 9129 6285 9163
rect 6285 9129 6319 9163
rect 6319 9129 6328 9163
rect 6276 9120 6328 9129
rect 8944 9120 8996 9172
rect 11704 9120 11756 9172
rect 4804 8984 4856 9036
rect 5632 8984 5684 9036
rect 10600 8984 10652 9036
rect 12808 9120 12860 9172
rect 16580 9120 16632 9172
rect 12624 9052 12676 9104
rect 12992 9052 13044 9104
rect 18236 9120 18288 9172
rect 23388 9163 23440 9172
rect 23388 9129 23397 9163
rect 23397 9129 23431 9163
rect 23431 9129 23440 9163
rect 23388 9120 23440 9129
rect 25136 9163 25188 9172
rect 25136 9129 25145 9163
rect 25145 9129 25179 9163
rect 25179 9129 25188 9163
rect 25136 9120 25188 9129
rect 5356 8916 5408 8968
rect 5816 8959 5868 8968
rect 5816 8925 5825 8959
rect 5825 8925 5859 8959
rect 5859 8925 5868 8959
rect 5816 8916 5868 8925
rect 5908 8959 5960 8968
rect 5908 8925 5917 8959
rect 5917 8925 5951 8959
rect 5951 8925 5960 8959
rect 5908 8916 5960 8925
rect 6092 8959 6144 8968
rect 6092 8925 6101 8959
rect 6101 8925 6135 8959
rect 6135 8925 6144 8959
rect 6092 8916 6144 8925
rect 8116 8959 8168 8968
rect 8116 8925 8125 8959
rect 8125 8925 8159 8959
rect 8159 8925 8168 8959
rect 8116 8916 8168 8925
rect 6184 8848 6236 8900
rect 8024 8848 8076 8900
rect 9680 8959 9732 8968
rect 9680 8925 9689 8959
rect 9689 8925 9723 8959
rect 9723 8925 9732 8959
rect 9680 8916 9732 8925
rect 9588 8848 9640 8900
rect 12072 8959 12124 8968
rect 12072 8925 12081 8959
rect 12081 8925 12115 8959
rect 12115 8925 12124 8959
rect 12072 8916 12124 8925
rect 12256 8959 12308 8968
rect 12256 8925 12265 8959
rect 12265 8925 12299 8959
rect 12299 8925 12308 8959
rect 12256 8916 12308 8925
rect 12348 8959 12400 8968
rect 12348 8925 12357 8959
rect 12357 8925 12391 8959
rect 12391 8925 12400 8959
rect 12348 8916 12400 8925
rect 13084 8959 13136 8968
rect 13084 8925 13093 8959
rect 13093 8925 13127 8959
rect 13127 8925 13136 8959
rect 13084 8916 13136 8925
rect 14096 8916 14148 8968
rect 17316 9052 17368 9104
rect 16580 8984 16632 9036
rect 16212 8916 16264 8968
rect 23388 8984 23440 9036
rect 24768 9027 24820 9036
rect 24768 8993 24777 9027
rect 24777 8993 24811 9027
rect 24811 8993 24820 9027
rect 24768 8984 24820 8993
rect 5908 8780 5960 8832
rect 11704 8780 11756 8832
rect 12440 8780 12492 8832
rect 17960 8848 18012 8900
rect 23664 8959 23716 8968
rect 23664 8925 23673 8959
rect 23673 8925 23707 8959
rect 23707 8925 23716 8959
rect 23664 8916 23716 8925
rect 23756 8891 23808 8900
rect 23756 8857 23765 8891
rect 23765 8857 23799 8891
rect 23799 8857 23808 8891
rect 23756 8848 23808 8857
rect 24032 8959 24084 8968
rect 24032 8925 24041 8959
rect 24041 8925 24075 8959
rect 24075 8925 24084 8959
rect 24032 8916 24084 8925
rect 24216 8959 24268 8968
rect 24216 8925 24225 8959
rect 24225 8925 24259 8959
rect 24259 8925 24268 8959
rect 24216 8916 24268 8925
rect 24124 8848 24176 8900
rect 17132 8780 17184 8832
rect 17592 8780 17644 8832
rect 18420 8780 18472 8832
rect 18788 8780 18840 8832
rect 23940 8780 23992 8832
rect 24216 8780 24268 8832
rect 24860 8959 24912 8968
rect 24860 8925 24869 8959
rect 24869 8925 24903 8959
rect 24903 8925 24912 8959
rect 24860 8916 24912 8925
rect 24952 8780 25004 8832
rect 4874 8678 4926 8730
rect 4938 8678 4990 8730
rect 5002 8678 5054 8730
rect 5066 8678 5118 8730
rect 5130 8678 5182 8730
rect 5816 8576 5868 8628
rect 9680 8619 9732 8628
rect 9680 8585 9689 8619
rect 9689 8585 9723 8619
rect 9723 8585 9732 8619
rect 9680 8576 9732 8585
rect 11704 8619 11756 8628
rect 11704 8585 11713 8619
rect 11713 8585 11747 8619
rect 11747 8585 11756 8619
rect 11704 8576 11756 8585
rect 14372 8576 14424 8628
rect 4804 8440 4856 8492
rect 5356 8483 5408 8492
rect 5356 8449 5365 8483
rect 5365 8449 5399 8483
rect 5399 8449 5408 8483
rect 5356 8440 5408 8449
rect 5540 8483 5592 8492
rect 5540 8449 5549 8483
rect 5549 8449 5583 8483
rect 5583 8449 5592 8483
rect 5540 8440 5592 8449
rect 5816 8440 5868 8492
rect 6000 8483 6052 8492
rect 6000 8449 6009 8483
rect 6009 8449 6043 8483
rect 6043 8449 6052 8483
rect 6000 8440 6052 8449
rect 6184 8483 6236 8492
rect 6184 8449 6193 8483
rect 6193 8449 6227 8483
rect 6227 8449 6236 8483
rect 6184 8440 6236 8449
rect 8024 8483 8076 8492
rect 8024 8449 8033 8483
rect 8033 8449 8067 8483
rect 8067 8449 8076 8483
rect 8024 8440 8076 8449
rect 5908 8372 5960 8424
rect 8116 8372 8168 8424
rect 9588 8508 9640 8560
rect 13084 8508 13136 8560
rect 9956 8483 10008 8492
rect 9956 8449 9965 8483
rect 9965 8449 9999 8483
rect 9999 8449 10008 8483
rect 9956 8440 10008 8449
rect 9588 8372 9640 8424
rect 12808 8483 12860 8492
rect 12808 8449 12817 8483
rect 12817 8449 12851 8483
rect 12851 8449 12860 8483
rect 12808 8440 12860 8449
rect 13912 8440 13964 8492
rect 24216 8576 24268 8628
rect 24860 8576 24912 8628
rect 17316 8551 17368 8560
rect 17316 8517 17325 8551
rect 17325 8517 17359 8551
rect 17359 8517 17368 8551
rect 17316 8508 17368 8517
rect 13820 8372 13872 8424
rect 14924 8440 14976 8492
rect 16856 8440 16908 8492
rect 9956 8304 10008 8356
rect 5816 8236 5868 8288
rect 10876 8236 10928 8288
rect 13452 8304 13504 8356
rect 13728 8304 13780 8356
rect 14924 8304 14976 8356
rect 17132 8483 17184 8492
rect 17132 8449 17141 8483
rect 17141 8449 17175 8483
rect 17175 8449 17184 8483
rect 17132 8440 17184 8449
rect 18972 8483 19024 8492
rect 18972 8449 18981 8483
rect 18981 8449 19015 8483
rect 19015 8449 19024 8483
rect 19984 8508 20036 8560
rect 18972 8440 19024 8449
rect 18144 8372 18196 8424
rect 18512 8372 18564 8424
rect 20904 8440 20956 8492
rect 23388 8551 23440 8560
rect 23388 8517 23397 8551
rect 23397 8517 23431 8551
rect 23431 8517 23440 8551
rect 23388 8508 23440 8517
rect 23940 8551 23992 8560
rect 23940 8517 23949 8551
rect 23949 8517 23983 8551
rect 23983 8517 23992 8551
rect 23940 8508 23992 8517
rect 20260 8372 20312 8424
rect 22008 8372 22060 8424
rect 23296 8483 23348 8492
rect 23296 8449 23305 8483
rect 23305 8449 23339 8483
rect 23339 8449 23348 8483
rect 23296 8440 23348 8449
rect 23572 8440 23624 8492
rect 25044 8440 25096 8492
rect 15936 8236 15988 8288
rect 16120 8236 16172 8288
rect 16764 8236 16816 8288
rect 19432 8304 19484 8356
rect 19708 8304 19760 8356
rect 20168 8304 20220 8356
rect 19524 8236 19576 8288
rect 19892 8279 19944 8288
rect 19892 8245 19901 8279
rect 19901 8245 19935 8279
rect 19935 8245 19944 8279
rect 19892 8236 19944 8245
rect 20628 8236 20680 8288
rect 20996 8236 21048 8288
rect 21180 8236 21232 8288
rect 22928 8304 22980 8356
rect 22284 8236 22336 8288
rect 23480 8304 23532 8356
rect 24032 8372 24084 8424
rect 24308 8236 24360 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 5356 8032 5408 8084
rect 6552 8032 6604 8084
rect 8484 8032 8536 8084
rect 9588 8032 9640 8084
rect 12624 8032 12676 8084
rect 13176 8075 13228 8084
rect 13176 8041 13185 8075
rect 13185 8041 13219 8075
rect 13219 8041 13228 8075
rect 13176 8032 13228 8041
rect 13912 8032 13964 8084
rect 17224 8075 17276 8084
rect 17224 8041 17233 8075
rect 17233 8041 17267 8075
rect 17267 8041 17276 8075
rect 17224 8032 17276 8041
rect 19892 8032 19944 8084
rect 20076 8075 20128 8084
rect 20076 8041 20085 8075
rect 20085 8041 20119 8075
rect 20119 8041 20128 8075
rect 20076 8032 20128 8041
rect 4620 7896 4672 7948
rect 16028 7964 16080 8016
rect 16948 7964 17000 8016
rect 4804 7871 4856 7880
rect 4804 7837 4813 7871
rect 4813 7837 4847 7871
rect 4847 7837 4856 7871
rect 4804 7828 4856 7837
rect 5816 7896 5868 7948
rect 5448 7871 5500 7880
rect 5448 7837 5457 7871
rect 5457 7837 5491 7871
rect 5491 7837 5500 7871
rect 5448 7828 5500 7837
rect 6092 7828 6144 7880
rect 9128 7828 9180 7880
rect 9588 7871 9640 7880
rect 9588 7837 9597 7871
rect 9597 7837 9631 7871
rect 9631 7837 9640 7871
rect 9588 7828 9640 7837
rect 12532 7871 12584 7880
rect 12532 7837 12541 7871
rect 12541 7837 12575 7871
rect 12575 7837 12584 7871
rect 12532 7828 12584 7837
rect 17684 7896 17736 7948
rect 12716 7871 12768 7880
rect 12716 7837 12725 7871
rect 12725 7837 12759 7871
rect 12759 7837 12768 7871
rect 12716 7828 12768 7837
rect 12900 7871 12952 7880
rect 12900 7837 12909 7871
rect 12909 7837 12943 7871
rect 12943 7837 12952 7871
rect 12900 7828 12952 7837
rect 12992 7871 13044 7880
rect 12992 7837 13001 7871
rect 13001 7837 13035 7871
rect 13035 7837 13044 7871
rect 12992 7828 13044 7837
rect 13820 7828 13872 7880
rect 15752 7871 15804 7880
rect 15752 7837 15761 7871
rect 15761 7837 15795 7871
rect 15795 7837 15804 7871
rect 15752 7828 15804 7837
rect 15936 7828 15988 7880
rect 16948 7828 17000 7880
rect 17040 7871 17092 7880
rect 17040 7837 17049 7871
rect 17049 7837 17083 7871
rect 17083 7837 17092 7871
rect 17040 7828 17092 7837
rect 17132 7828 17184 7880
rect 17592 7871 17644 7880
rect 17592 7837 17601 7871
rect 17601 7837 17635 7871
rect 17635 7837 17644 7871
rect 17592 7828 17644 7837
rect 17776 7871 17828 7880
rect 17776 7837 17785 7871
rect 17785 7837 17819 7871
rect 17819 7837 17828 7871
rect 17776 7828 17828 7837
rect 9956 7692 10008 7744
rect 10600 7692 10652 7744
rect 12348 7760 12400 7812
rect 13728 7803 13780 7812
rect 13728 7769 13737 7803
rect 13737 7769 13771 7803
rect 13771 7769 13780 7803
rect 13728 7760 13780 7769
rect 13176 7692 13228 7744
rect 13360 7735 13412 7744
rect 13360 7701 13369 7735
rect 13369 7701 13403 7735
rect 13403 7701 13412 7735
rect 13360 7692 13412 7701
rect 14188 7760 14240 7812
rect 16580 7760 16632 7812
rect 18420 7871 18472 7880
rect 18420 7837 18429 7871
rect 18429 7837 18463 7871
rect 18463 7837 18472 7871
rect 18420 7828 18472 7837
rect 18512 7871 18564 7880
rect 18512 7837 18521 7871
rect 18521 7837 18555 7871
rect 18555 7837 18564 7871
rect 18512 7828 18564 7837
rect 18604 7871 18656 7880
rect 18604 7837 18613 7871
rect 18613 7837 18647 7871
rect 18647 7837 18656 7871
rect 18604 7828 18656 7837
rect 18788 7871 18840 7880
rect 18788 7837 18797 7871
rect 18797 7837 18831 7871
rect 18831 7837 18840 7871
rect 18788 7828 18840 7837
rect 18880 7871 18932 7880
rect 18880 7837 18889 7871
rect 18889 7837 18923 7871
rect 18923 7837 18932 7871
rect 18880 7828 18932 7837
rect 18052 7760 18104 7812
rect 18236 7760 18288 7812
rect 19156 7760 19208 7812
rect 14556 7692 14608 7744
rect 15200 7692 15252 7744
rect 15936 7692 15988 7744
rect 16672 7692 16724 7744
rect 17040 7692 17092 7744
rect 17408 7692 17460 7744
rect 19064 7735 19116 7744
rect 19064 7701 19073 7735
rect 19073 7701 19107 7735
rect 19107 7701 19116 7735
rect 19064 7692 19116 7701
rect 19248 7735 19300 7744
rect 19248 7701 19257 7735
rect 19257 7701 19291 7735
rect 19291 7701 19300 7735
rect 19248 7692 19300 7701
rect 22192 8075 22244 8084
rect 22192 8041 22201 8075
rect 22201 8041 22235 8075
rect 22235 8041 22244 8075
rect 22192 8032 22244 8041
rect 21272 7964 21324 8016
rect 19708 7939 19760 7948
rect 19708 7905 19717 7939
rect 19717 7905 19751 7939
rect 19751 7905 19760 7939
rect 19708 7896 19760 7905
rect 21180 7896 21232 7948
rect 19524 7871 19576 7880
rect 19524 7837 19533 7871
rect 19533 7837 19567 7871
rect 19567 7837 19576 7871
rect 19524 7828 19576 7837
rect 19616 7828 19668 7880
rect 19984 7871 20036 7880
rect 19984 7837 19993 7871
rect 19993 7837 20027 7871
rect 20027 7837 20036 7871
rect 19984 7828 20036 7837
rect 19432 7760 19484 7812
rect 20444 7828 20496 7880
rect 20536 7871 20588 7880
rect 20536 7837 20545 7871
rect 20545 7837 20579 7871
rect 20579 7837 20588 7871
rect 20536 7828 20588 7837
rect 20628 7871 20680 7880
rect 20628 7837 20637 7871
rect 20637 7837 20671 7871
rect 20671 7837 20680 7871
rect 20628 7828 20680 7837
rect 21088 7828 21140 7880
rect 21548 7828 21600 7880
rect 23388 7964 23440 8016
rect 23756 8075 23808 8084
rect 23756 8041 23765 8075
rect 23765 8041 23799 8075
rect 23799 8041 23808 8075
rect 23756 8032 23808 8041
rect 25044 8032 25096 8084
rect 23848 7964 23900 8016
rect 24308 7964 24360 8016
rect 23480 7896 23532 7948
rect 24768 7896 24820 7948
rect 23756 7828 23808 7880
rect 24124 7871 24176 7880
rect 24124 7837 24133 7871
rect 24133 7837 24167 7871
rect 24167 7837 24176 7871
rect 24124 7828 24176 7837
rect 25688 7828 25740 7880
rect 27712 7828 27764 7880
rect 21640 7760 21692 7812
rect 23296 7760 23348 7812
rect 27620 7760 27672 7812
rect 21732 7692 21784 7744
rect 22744 7735 22796 7744
rect 22744 7701 22753 7735
rect 22753 7701 22787 7735
rect 22787 7701 22796 7735
rect 22744 7692 22796 7701
rect 23756 7692 23808 7744
rect 4874 7590 4926 7642
rect 4938 7590 4990 7642
rect 5002 7590 5054 7642
rect 5066 7590 5118 7642
rect 5130 7590 5182 7642
rect 4804 7488 4856 7540
rect 5264 7488 5316 7540
rect 8024 7488 8076 7540
rect 8300 7531 8352 7540
rect 8300 7497 8309 7531
rect 8309 7497 8343 7531
rect 8343 7497 8352 7531
rect 8852 7531 8904 7540
rect 8300 7488 8352 7497
rect 8852 7497 8861 7531
rect 8861 7497 8895 7531
rect 8895 7497 8904 7531
rect 8852 7488 8904 7497
rect 5540 7352 5592 7404
rect 5448 7284 5500 7336
rect 5816 7352 5868 7404
rect 6552 7395 6604 7404
rect 6552 7361 6561 7395
rect 6561 7361 6595 7395
rect 6595 7361 6604 7395
rect 6552 7352 6604 7361
rect 5540 7148 5592 7200
rect 7564 7216 7616 7268
rect 8024 7352 8076 7404
rect 8392 7395 8444 7404
rect 8392 7361 8401 7395
rect 8401 7361 8435 7395
rect 8435 7361 8444 7395
rect 8392 7352 8444 7361
rect 8484 7395 8536 7404
rect 8484 7361 8493 7395
rect 8493 7361 8527 7395
rect 8527 7361 8536 7395
rect 8484 7352 8536 7361
rect 8576 7352 8628 7404
rect 9036 7352 9088 7404
rect 9128 7395 9180 7404
rect 9128 7361 9137 7395
rect 9137 7361 9171 7395
rect 9171 7361 9180 7395
rect 9128 7352 9180 7361
rect 9772 7488 9824 7540
rect 12164 7531 12216 7540
rect 12164 7497 12173 7531
rect 12173 7497 12207 7531
rect 12207 7497 12216 7531
rect 12164 7488 12216 7497
rect 12992 7488 13044 7540
rect 14096 7531 14148 7540
rect 14096 7497 14105 7531
rect 14105 7497 14139 7531
rect 14139 7497 14148 7531
rect 14096 7488 14148 7497
rect 14556 7531 14608 7540
rect 14556 7497 14565 7531
rect 14565 7497 14599 7531
rect 14599 7497 14608 7531
rect 14556 7488 14608 7497
rect 15016 7488 15068 7540
rect 16212 7488 16264 7540
rect 17684 7488 17736 7540
rect 18052 7531 18104 7540
rect 18052 7497 18061 7531
rect 18061 7497 18095 7531
rect 18095 7497 18104 7531
rect 18052 7488 18104 7497
rect 18144 7488 18196 7540
rect 18420 7488 18472 7540
rect 20076 7488 20128 7540
rect 20536 7488 20588 7540
rect 10600 7463 10652 7472
rect 10600 7429 10609 7463
rect 10609 7429 10643 7463
rect 10643 7429 10652 7463
rect 10600 7420 10652 7429
rect 10876 7420 10928 7472
rect 12440 7420 12492 7472
rect 9680 7395 9732 7404
rect 9680 7361 9689 7395
rect 9689 7361 9723 7395
rect 9723 7361 9732 7395
rect 9680 7352 9732 7361
rect 9588 7284 9640 7336
rect 10692 7352 10744 7404
rect 11612 7395 11664 7404
rect 11612 7361 11621 7395
rect 11621 7361 11655 7395
rect 11655 7361 11664 7395
rect 11612 7352 11664 7361
rect 11888 7395 11940 7404
rect 11888 7361 11897 7395
rect 11897 7361 11931 7395
rect 11931 7361 11940 7395
rect 11888 7352 11940 7361
rect 13084 7420 13136 7472
rect 13360 7352 13412 7404
rect 13452 7395 13504 7404
rect 13452 7361 13461 7395
rect 13461 7361 13495 7395
rect 13495 7361 13504 7395
rect 13452 7352 13504 7361
rect 11704 7284 11756 7336
rect 13820 7395 13872 7404
rect 13820 7361 13829 7395
rect 13829 7361 13863 7395
rect 13863 7361 13872 7395
rect 13820 7352 13872 7361
rect 13912 7395 13964 7404
rect 13912 7361 13921 7395
rect 13921 7361 13955 7395
rect 13955 7361 13964 7395
rect 13912 7352 13964 7361
rect 14556 7352 14608 7404
rect 13728 7284 13780 7336
rect 14740 7420 14792 7472
rect 14832 7395 14884 7404
rect 14832 7361 14841 7395
rect 14841 7361 14875 7395
rect 14875 7361 14884 7395
rect 14832 7352 14884 7361
rect 15200 7463 15252 7472
rect 15200 7429 15209 7463
rect 15209 7429 15243 7463
rect 15243 7429 15252 7463
rect 15200 7420 15252 7429
rect 15108 7395 15160 7404
rect 15108 7361 15117 7395
rect 15117 7361 15151 7395
rect 15151 7361 15160 7395
rect 15108 7352 15160 7361
rect 15384 7352 15436 7404
rect 15568 7395 15620 7404
rect 15568 7361 15577 7395
rect 15577 7361 15611 7395
rect 15611 7361 15620 7395
rect 15568 7352 15620 7361
rect 15844 7395 15896 7404
rect 15844 7361 15853 7395
rect 15853 7361 15887 7395
rect 15887 7361 15896 7395
rect 15844 7352 15896 7361
rect 15936 7395 15988 7404
rect 15936 7361 15945 7395
rect 15945 7361 15979 7395
rect 15979 7361 15988 7395
rect 15936 7352 15988 7361
rect 16212 7395 16264 7404
rect 16212 7361 16221 7395
rect 16221 7361 16255 7395
rect 16255 7361 16264 7395
rect 16212 7352 16264 7361
rect 16580 7352 16632 7404
rect 16764 7395 16816 7404
rect 16764 7361 16773 7395
rect 16773 7361 16807 7395
rect 16807 7361 16816 7395
rect 16764 7352 16816 7361
rect 17040 7352 17092 7404
rect 17408 7352 17460 7404
rect 6552 7148 6604 7200
rect 9036 7148 9088 7200
rect 14372 7216 14424 7268
rect 16856 7216 16908 7268
rect 17040 7216 17092 7268
rect 17316 7327 17368 7336
rect 17316 7293 17325 7327
rect 17325 7293 17359 7327
rect 17359 7293 17368 7327
rect 17316 7284 17368 7293
rect 12440 7148 12492 7200
rect 12992 7148 13044 7200
rect 13084 7191 13136 7200
rect 13084 7157 13093 7191
rect 13093 7157 13127 7191
rect 13127 7157 13136 7191
rect 13084 7148 13136 7157
rect 13268 7191 13320 7200
rect 13268 7157 13277 7191
rect 13277 7157 13311 7191
rect 13311 7157 13320 7191
rect 13268 7148 13320 7157
rect 16028 7148 16080 7200
rect 16304 7148 16356 7200
rect 18512 7420 18564 7472
rect 17592 7395 17644 7404
rect 17592 7361 17601 7395
rect 17601 7361 17635 7395
rect 17635 7361 17644 7395
rect 17592 7352 17644 7361
rect 17868 7352 17920 7404
rect 17960 7352 18012 7404
rect 18236 7395 18288 7404
rect 18236 7361 18245 7395
rect 18245 7361 18279 7395
rect 18279 7361 18288 7395
rect 18236 7352 18288 7361
rect 19064 7395 19116 7404
rect 19064 7361 19073 7395
rect 19073 7361 19107 7395
rect 19107 7361 19116 7395
rect 19064 7352 19116 7361
rect 23296 7531 23348 7540
rect 23296 7497 23305 7531
rect 23305 7497 23339 7531
rect 23339 7497 23348 7531
rect 23296 7488 23348 7497
rect 24768 7488 24820 7540
rect 21180 7420 21232 7472
rect 18604 7284 18656 7336
rect 19248 7327 19300 7336
rect 19248 7293 19257 7327
rect 19257 7293 19291 7327
rect 19291 7293 19300 7327
rect 19248 7284 19300 7293
rect 19800 7284 19852 7336
rect 20812 7395 20864 7404
rect 20812 7361 20821 7395
rect 20821 7361 20855 7395
rect 20855 7361 20864 7395
rect 20812 7352 20864 7361
rect 20904 7352 20956 7404
rect 21088 7395 21140 7404
rect 21088 7361 21097 7395
rect 21097 7361 21131 7395
rect 21131 7361 21140 7395
rect 21088 7352 21140 7361
rect 20536 7284 20588 7336
rect 20444 7216 20496 7268
rect 21640 7395 21692 7404
rect 21640 7361 21649 7395
rect 21649 7361 21683 7395
rect 21683 7361 21692 7395
rect 21640 7352 21692 7361
rect 22008 7395 22060 7404
rect 22008 7361 22017 7395
rect 22017 7361 22051 7395
rect 22051 7361 22060 7395
rect 22008 7352 22060 7361
rect 23756 7463 23808 7472
rect 23756 7429 23765 7463
rect 23765 7429 23799 7463
rect 23799 7429 23808 7463
rect 23756 7420 23808 7429
rect 25044 7420 25096 7472
rect 22284 7395 22336 7404
rect 22284 7361 22293 7395
rect 22293 7361 22327 7395
rect 22327 7361 22336 7395
rect 22284 7352 22336 7361
rect 22468 7395 22520 7404
rect 22468 7361 22477 7395
rect 22477 7361 22511 7395
rect 22511 7361 22520 7395
rect 22468 7352 22520 7361
rect 23388 7395 23440 7404
rect 23388 7361 23397 7395
rect 23397 7361 23431 7395
rect 23431 7361 23440 7395
rect 23388 7352 23440 7361
rect 23480 7395 23532 7404
rect 23480 7361 23489 7395
rect 23489 7361 23523 7395
rect 23523 7361 23532 7395
rect 23480 7352 23532 7361
rect 21732 7284 21784 7336
rect 22376 7216 22428 7268
rect 21180 7148 21232 7200
rect 21364 7191 21416 7200
rect 21364 7157 21373 7191
rect 21373 7157 21407 7191
rect 21407 7157 21416 7191
rect 21364 7148 21416 7157
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 8024 6987 8076 6996
rect 8024 6953 8033 6987
rect 8033 6953 8067 6987
rect 8067 6953 8076 6987
rect 8024 6944 8076 6953
rect 9128 6944 9180 6996
rect 9588 6944 9640 6996
rect 5264 6876 5316 6928
rect 5540 6851 5592 6860
rect 5540 6817 5549 6851
rect 5549 6817 5583 6851
rect 5583 6817 5592 6851
rect 5540 6808 5592 6817
rect 7564 6876 7616 6928
rect 8484 6876 8536 6928
rect 7564 6783 7616 6792
rect 7564 6749 7573 6783
rect 7573 6749 7607 6783
rect 7607 6749 7616 6783
rect 7564 6740 7616 6749
rect 8392 6808 8444 6860
rect 11888 6919 11940 6928
rect 11888 6885 11897 6919
rect 11897 6885 11931 6919
rect 11931 6885 11940 6919
rect 11888 6876 11940 6885
rect 12900 6944 12952 6996
rect 13084 6944 13136 6996
rect 15016 6987 15068 6996
rect 15016 6953 15025 6987
rect 15025 6953 15059 6987
rect 15059 6953 15068 6987
rect 15016 6944 15068 6953
rect 15108 6944 15160 6996
rect 15384 6944 15436 6996
rect 15752 6944 15804 6996
rect 16672 6944 16724 6996
rect 17316 6944 17368 6996
rect 17592 6944 17644 6996
rect 21364 6944 21416 6996
rect 21548 6944 21600 6996
rect 22468 6944 22520 6996
rect 12256 6876 12308 6928
rect 8576 6783 8628 6792
rect 8576 6749 8585 6783
rect 8585 6749 8619 6783
rect 8619 6749 8628 6783
rect 8576 6740 8628 6749
rect 8760 6783 8812 6792
rect 8760 6749 8769 6783
rect 8769 6749 8803 6783
rect 8803 6749 8812 6783
rect 8760 6740 8812 6749
rect 8852 6740 8904 6792
rect 9680 6740 9732 6792
rect 9772 6783 9824 6792
rect 9772 6749 9781 6783
rect 9781 6749 9815 6783
rect 9815 6749 9824 6783
rect 9772 6740 9824 6749
rect 10324 6783 10376 6792
rect 10324 6749 10333 6783
rect 10333 6749 10367 6783
rect 10367 6749 10376 6783
rect 10324 6740 10376 6749
rect 12440 6740 12492 6792
rect 12624 6876 12676 6928
rect 14372 6876 14424 6928
rect 15568 6876 15620 6928
rect 15844 6876 15896 6928
rect 14188 6851 14240 6860
rect 12900 6783 12952 6792
rect 12900 6749 12909 6783
rect 12909 6749 12943 6783
rect 12943 6749 12952 6783
rect 12900 6740 12952 6749
rect 12992 6783 13044 6792
rect 12992 6749 13001 6783
rect 13001 6749 13035 6783
rect 13035 6749 13044 6783
rect 12992 6740 13044 6749
rect 13268 6783 13320 6792
rect 13268 6749 13277 6783
rect 13277 6749 13311 6783
rect 13311 6749 13320 6783
rect 13268 6740 13320 6749
rect 8484 6715 8536 6724
rect 8484 6681 8493 6715
rect 8493 6681 8527 6715
rect 8527 6681 8536 6715
rect 8484 6672 8536 6681
rect 13452 6715 13504 6724
rect 6000 6647 6052 6656
rect 6000 6613 6009 6647
rect 6009 6613 6043 6647
rect 6043 6613 6052 6647
rect 6000 6604 6052 6613
rect 8392 6604 8444 6656
rect 8668 6647 8720 6656
rect 8668 6613 8677 6647
rect 8677 6613 8711 6647
rect 8711 6613 8720 6647
rect 8668 6604 8720 6613
rect 10232 6647 10284 6656
rect 10232 6613 10241 6647
rect 10241 6613 10275 6647
rect 10275 6613 10284 6647
rect 10232 6604 10284 6613
rect 13452 6681 13461 6715
rect 13461 6681 13495 6715
rect 13495 6681 13504 6715
rect 13452 6672 13504 6681
rect 12716 6604 12768 6656
rect 13728 6740 13780 6792
rect 14188 6817 14197 6851
rect 14197 6817 14231 6851
rect 14231 6817 14240 6851
rect 14188 6808 14240 6817
rect 14280 6783 14332 6792
rect 14280 6749 14289 6783
rect 14289 6749 14323 6783
rect 14323 6749 14332 6783
rect 14280 6740 14332 6749
rect 14924 6783 14976 6792
rect 14924 6749 14933 6783
rect 14933 6749 14967 6783
rect 14967 6749 14976 6783
rect 14924 6740 14976 6749
rect 18144 6808 18196 6860
rect 18972 6808 19024 6860
rect 20352 6808 20404 6860
rect 15476 6783 15528 6792
rect 15476 6749 15485 6783
rect 15485 6749 15519 6783
rect 15519 6749 15528 6783
rect 15476 6740 15528 6749
rect 15844 6783 15896 6792
rect 15844 6749 15853 6783
rect 15853 6749 15887 6783
rect 15887 6749 15896 6783
rect 15844 6740 15896 6749
rect 16488 6740 16540 6792
rect 18696 6740 18748 6792
rect 21456 6740 21508 6792
rect 23388 6740 23440 6792
rect 24308 6740 24360 6792
rect 16212 6672 16264 6724
rect 16304 6604 16356 6656
rect 4874 6502 4926 6554
rect 4938 6502 4990 6554
rect 5002 6502 5054 6554
rect 5066 6502 5118 6554
rect 5130 6502 5182 6554
rect 6000 6264 6052 6316
rect 8576 6264 8628 6316
rect 8944 6307 8996 6316
rect 8944 6273 8953 6307
rect 8953 6273 8987 6307
rect 8987 6273 8996 6307
rect 8944 6264 8996 6273
rect 10232 6264 10284 6316
rect 12532 6400 12584 6452
rect 11888 6332 11940 6384
rect 13176 6332 13228 6384
rect 13452 6307 13504 6316
rect 13452 6273 13461 6307
rect 13461 6273 13495 6307
rect 13495 6273 13504 6307
rect 13452 6264 13504 6273
rect 8392 6239 8444 6248
rect 8392 6205 8401 6239
rect 8401 6205 8435 6239
rect 8435 6205 8444 6239
rect 8392 6196 8444 6205
rect 9680 6196 9732 6248
rect 10324 6196 10376 6248
rect 8760 6128 8812 6180
rect 13728 6264 13780 6316
rect 14280 6196 14332 6248
rect 16028 6375 16080 6384
rect 16028 6341 16037 6375
rect 16037 6341 16071 6375
rect 16071 6341 16080 6375
rect 16028 6332 16080 6341
rect 18604 6443 18656 6452
rect 18604 6409 18613 6443
rect 18613 6409 18647 6443
rect 18647 6409 18656 6443
rect 18604 6400 18656 6409
rect 27620 6443 27672 6452
rect 27620 6409 27629 6443
rect 27629 6409 27663 6443
rect 27663 6409 27672 6443
rect 27620 6400 27672 6409
rect 17040 6332 17092 6384
rect 16488 6264 16540 6316
rect 18696 6332 18748 6384
rect 27804 6307 27856 6316
rect 27804 6273 27813 6307
rect 27813 6273 27847 6307
rect 27847 6273 27856 6307
rect 27804 6264 27856 6273
rect 13820 6128 13872 6180
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 8484 5856 8536 5908
rect 13268 5856 13320 5908
rect 15476 5856 15528 5908
rect 27712 5856 27764 5908
rect 8392 5695 8444 5704
rect 8392 5661 8401 5695
rect 8401 5661 8435 5695
rect 8435 5661 8444 5695
rect 8392 5652 8444 5661
rect 8944 5720 8996 5772
rect 8668 5695 8720 5704
rect 8668 5661 8677 5695
rect 8677 5661 8711 5695
rect 8711 5661 8720 5695
rect 8668 5652 8720 5661
rect 27804 5695 27856 5704
rect 27804 5661 27813 5695
rect 27813 5661 27847 5695
rect 27847 5661 27856 5695
rect 27804 5652 27856 5661
rect 4874 5414 4926 5466
rect 4938 5414 4990 5466
rect 5002 5414 5054 5466
rect 5066 5414 5118 5466
rect 5130 5414 5182 5466
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 4874 4326 4926 4378
rect 4938 4326 4990 4378
rect 5002 4326 5054 4378
rect 5066 4326 5118 4378
rect 5130 4326 5182 4378
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 4874 3238 4926 3290
rect 4938 3238 4990 3290
rect 5002 3238 5054 3290
rect 5066 3238 5118 3290
rect 5130 3238 5182 3290
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 6092 2635 6144 2644
rect 6092 2601 6101 2635
rect 6101 2601 6135 2635
rect 6135 2601 6144 2635
rect 6092 2592 6144 2601
rect 9312 2635 9364 2644
rect 9312 2601 9321 2635
rect 9321 2601 9355 2635
rect 9355 2601 9364 2635
rect 9312 2592 9364 2601
rect 5816 2388 5868 2440
rect 9036 2388 9088 2440
rect 4874 2150 4926 2202
rect 4938 2150 4990 2202
rect 5002 2150 5054 2202
rect 5066 2150 5118 2202
rect 5130 2150 5182 2202
<< metal2 >>
rect 11610 30818 11666 31476
rect 12254 30818 12310 31476
rect 12898 30818 12954 31476
rect 13542 30818 13598 31476
rect 14186 30818 14242 31476
rect 14830 30818 14886 31476
rect 15474 30818 15530 31476
rect 16118 30818 16174 31476
rect 16762 30818 16818 31476
rect 17406 30818 17462 31476
rect 18050 30818 18106 31476
rect 18694 30818 18750 31476
rect 19338 30818 19394 31476
rect 19982 30818 20038 31476
rect 20626 30818 20682 31476
rect 11610 30790 11836 30818
rect 11610 30676 11666 30790
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 11808 28762 11836 30790
rect 12254 30790 12388 30818
rect 12254 30676 12310 30790
rect 12360 28762 12388 30790
rect 12898 30790 13124 30818
rect 12898 30676 12954 30790
rect 13096 28762 13124 30790
rect 13542 30790 13768 30818
rect 13542 30676 13598 30790
rect 13740 28762 13768 30790
rect 14186 30790 14412 30818
rect 14186 30676 14242 30790
rect 14384 28762 14412 30790
rect 14830 30790 15056 30818
rect 14830 30676 14886 30790
rect 15028 28762 15056 30790
rect 15474 30790 15700 30818
rect 15474 30676 15530 30790
rect 15672 28762 15700 30790
rect 16118 30790 16344 30818
rect 16118 30676 16174 30790
rect 16316 28762 16344 30790
rect 16762 30790 16988 30818
rect 16762 30676 16818 30790
rect 16960 28762 16988 30790
rect 17406 30790 17632 30818
rect 17406 30676 17462 30790
rect 17604 28762 17632 30790
rect 18050 30790 18276 30818
rect 18050 30676 18106 30790
rect 18248 28762 18276 30790
rect 18694 30790 18920 30818
rect 18694 30676 18750 30790
rect 18892 28762 18920 30790
rect 19338 30790 19656 30818
rect 19338 30676 19394 30790
rect 19628 28762 19656 30790
rect 19982 30790 20300 30818
rect 19982 30676 20038 30790
rect 20272 28762 20300 30790
rect 20548 30790 20682 30818
rect 20548 28762 20576 30790
rect 20626 30676 20682 30790
rect 21270 30818 21326 31476
rect 21914 30818 21970 31476
rect 22558 30818 22614 31476
rect 23202 30818 23258 31476
rect 23846 30818 23902 31476
rect 24490 30818 24546 31476
rect 25134 30818 25190 31476
rect 25778 30818 25834 31476
rect 26422 30818 26478 31476
rect 27066 30818 27122 31476
rect 27710 30818 27766 31476
rect 28354 30818 28410 31476
rect 28998 30818 29054 31476
rect 21270 30790 21588 30818
rect 21270 30676 21326 30790
rect 21560 28762 21588 30790
rect 21914 30790 22048 30818
rect 21914 30676 21970 30790
rect 22020 28762 22048 30790
rect 22558 30790 22876 30818
rect 22558 30676 22614 30790
rect 22848 28762 22876 30790
rect 23202 30790 23428 30818
rect 23202 30676 23258 30790
rect 23400 28762 23428 30790
rect 23846 30790 24164 30818
rect 23846 30676 23902 30790
rect 24136 28762 24164 30790
rect 24490 30790 24808 30818
rect 24490 30676 24546 30790
rect 24780 28762 24808 30790
rect 25134 30790 25452 30818
rect 25134 30676 25190 30790
rect 25424 28762 25452 30790
rect 25778 30790 26096 30818
rect 25778 30676 25834 30790
rect 26068 28762 26096 30790
rect 26422 30790 26740 30818
rect 26422 30676 26478 30790
rect 26712 28762 26740 30790
rect 27066 30790 27384 30818
rect 27066 30676 27122 30790
rect 27356 28762 27384 30790
rect 27710 30790 27844 30818
rect 27710 30676 27766 30790
rect 27816 28762 27844 30790
rect 28000 30790 28410 30818
rect 11796 28756 11848 28762
rect 11796 28698 11848 28704
rect 12348 28756 12400 28762
rect 12348 28698 12400 28704
rect 13084 28756 13136 28762
rect 13084 28698 13136 28704
rect 13728 28756 13780 28762
rect 13728 28698 13780 28704
rect 14372 28756 14424 28762
rect 14372 28698 14424 28704
rect 15016 28756 15068 28762
rect 15016 28698 15068 28704
rect 15660 28756 15712 28762
rect 15660 28698 15712 28704
rect 16304 28756 16356 28762
rect 16304 28698 16356 28704
rect 16948 28756 17000 28762
rect 16948 28698 17000 28704
rect 17592 28756 17644 28762
rect 17592 28698 17644 28704
rect 18236 28756 18288 28762
rect 18236 28698 18288 28704
rect 18880 28756 18932 28762
rect 18880 28698 18932 28704
rect 19616 28756 19668 28762
rect 19616 28698 19668 28704
rect 20260 28756 20312 28762
rect 20260 28698 20312 28704
rect 20536 28756 20588 28762
rect 20536 28698 20588 28704
rect 21548 28756 21600 28762
rect 21548 28698 21600 28704
rect 22008 28756 22060 28762
rect 22008 28698 22060 28704
rect 22836 28756 22888 28762
rect 22836 28698 22888 28704
rect 23388 28756 23440 28762
rect 23388 28698 23440 28704
rect 24124 28756 24176 28762
rect 24124 28698 24176 28704
rect 24768 28756 24820 28762
rect 24768 28698 24820 28704
rect 25412 28756 25464 28762
rect 25412 28698 25464 28704
rect 26056 28756 26108 28762
rect 26056 28698 26108 28704
rect 26700 28756 26752 28762
rect 26700 28698 26752 28704
rect 27344 28756 27396 28762
rect 27344 28698 27396 28704
rect 27804 28756 27856 28762
rect 27804 28698 27856 28704
rect 18144 28688 18196 28694
rect 18144 28630 18196 28636
rect 17960 28620 18012 28626
rect 17960 28562 18012 28568
rect 11980 28552 12032 28558
rect 11980 28494 12032 28500
rect 13268 28552 13320 28558
rect 13268 28494 13320 28500
rect 15844 28552 15896 28558
rect 15844 28494 15896 28500
rect 16948 28552 17000 28558
rect 16948 28494 17000 28500
rect 17132 28552 17184 28558
rect 17132 28494 17184 28500
rect 17868 28552 17920 28558
rect 17868 28494 17920 28500
rect 4874 28316 5182 28325
rect 4874 28314 4880 28316
rect 4936 28314 4960 28316
rect 5016 28314 5040 28316
rect 5096 28314 5120 28316
rect 5176 28314 5182 28316
rect 4936 28262 4938 28314
rect 5118 28262 5120 28314
rect 4874 28260 4880 28262
rect 4936 28260 4960 28262
rect 5016 28260 5040 28262
rect 5096 28260 5120 28262
rect 5176 28260 5182 28262
rect 4874 28251 5182 28260
rect 11992 28082 12020 28494
rect 13280 28150 13308 28494
rect 13268 28144 13320 28150
rect 13268 28086 13320 28092
rect 11060 28076 11112 28082
rect 11060 28018 11112 28024
rect 11704 28076 11756 28082
rect 11704 28018 11756 28024
rect 11980 28076 12032 28082
rect 11980 28018 12032 28024
rect 7472 28008 7524 28014
rect 7472 27950 7524 27956
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 2780 27668 2832 27674
rect 2780 27610 2832 27616
rect 6920 27668 6972 27674
rect 6920 27610 6972 27616
rect 2044 27464 2096 27470
rect 2044 27406 2096 27412
rect 2056 26994 2084 27406
rect 2792 27062 2820 27610
rect 3148 27600 3200 27606
rect 5448 27600 5500 27606
rect 3148 27542 3200 27548
rect 5184 27560 5448 27588
rect 2780 27056 2832 27062
rect 2780 26998 2832 27004
rect 2044 26988 2096 26994
rect 2044 26930 2096 26936
rect 1768 26240 1820 26246
rect 1768 26182 1820 26188
rect 1780 24206 1808 26182
rect 848 24200 900 24206
rect 848 24142 900 24148
rect 1768 24200 1820 24206
rect 1768 24142 1820 24148
rect 860 24041 888 24142
rect 1584 24064 1636 24070
rect 846 24032 902 24041
rect 1584 24006 1636 24012
rect 846 23967 902 23976
rect 1596 23866 1624 24006
rect 1584 23860 1636 23866
rect 1584 23802 1636 23808
rect 1492 23724 1544 23730
rect 1492 23666 1544 23672
rect 1504 23225 1532 23666
rect 1490 23216 1546 23225
rect 1490 23151 1546 23160
rect 848 22704 900 22710
rect 846 22672 848 22681
rect 900 22672 902 22681
rect 846 22607 902 22616
rect 848 22024 900 22030
rect 846 21992 848 22001
rect 900 21992 902 22001
rect 846 21927 902 21936
rect 1030 21176 1086 21185
rect 1030 21111 1086 21120
rect 1044 20942 1072 21111
rect 1032 20936 1084 20942
rect 1032 20878 1084 20884
rect 1780 20874 1808 24142
rect 2056 23526 2084 26930
rect 2136 26920 2188 26926
rect 2136 26862 2188 26868
rect 2596 26920 2648 26926
rect 2596 26862 2648 26868
rect 2148 26518 2176 26862
rect 2504 26784 2556 26790
rect 2504 26726 2556 26732
rect 2136 26512 2188 26518
rect 2136 26454 2188 26460
rect 2044 23520 2096 23526
rect 2044 23462 2096 23468
rect 2056 21570 2084 23462
rect 2148 22438 2176 26454
rect 2516 26314 2544 26726
rect 2608 26518 2636 26862
rect 2596 26512 2648 26518
rect 2596 26454 2648 26460
rect 2504 26308 2556 26314
rect 2504 26250 2556 26256
rect 2516 25362 2544 26250
rect 2792 26246 2820 26998
rect 3056 26852 3108 26858
rect 3056 26794 3108 26800
rect 3068 26586 3096 26794
rect 3056 26580 3108 26586
rect 3056 26522 3108 26528
rect 2780 26240 2832 26246
rect 2780 26182 2832 26188
rect 2792 26042 2820 26182
rect 2780 26036 2832 26042
rect 2780 25978 2832 25984
rect 2504 25356 2556 25362
rect 2504 25298 2556 25304
rect 2792 25294 2820 25978
rect 2780 25288 2832 25294
rect 2780 25230 2832 25236
rect 2596 24200 2648 24206
rect 2596 24142 2648 24148
rect 3056 24200 3108 24206
rect 3056 24142 3108 24148
rect 2504 24132 2556 24138
rect 2504 24074 2556 24080
rect 2516 23730 2544 24074
rect 2504 23724 2556 23730
rect 2504 23666 2556 23672
rect 2228 22636 2280 22642
rect 2228 22578 2280 22584
rect 2136 22432 2188 22438
rect 2136 22374 2188 22380
rect 2240 22098 2268 22578
rect 2412 22432 2464 22438
rect 2412 22374 2464 22380
rect 2228 22092 2280 22098
rect 2228 22034 2280 22040
rect 2240 21690 2268 22034
rect 2228 21684 2280 21690
rect 2228 21626 2280 21632
rect 2056 21542 2268 21570
rect 1492 20868 1544 20874
rect 1492 20810 1544 20816
rect 1768 20868 1820 20874
rect 1768 20810 1820 20816
rect 2136 20868 2188 20874
rect 2136 20810 2188 20816
rect 1504 20505 1532 20810
rect 1952 20528 2004 20534
rect 1490 20496 1546 20505
rect 1952 20470 2004 20476
rect 1490 20431 1546 20440
rect 1584 19984 1636 19990
rect 846 19952 902 19961
rect 1584 19926 1636 19932
rect 846 19887 902 19896
rect 860 19854 888 19887
rect 848 19848 900 19854
rect 848 19790 900 19796
rect 1596 19514 1624 19926
rect 1964 19854 1992 20470
rect 1952 19848 2004 19854
rect 2004 19796 2084 19802
rect 1952 19790 2084 19796
rect 1964 19774 2084 19790
rect 1584 19508 1636 19514
rect 1584 19450 1636 19456
rect 1400 19372 1452 19378
rect 1400 19314 1452 19320
rect 1412 19145 1440 19314
rect 1398 19136 1454 19145
rect 1398 19071 1454 19080
rect 1596 17678 1624 19450
rect 2056 19310 2084 19774
rect 2044 19304 2096 19310
rect 2044 19246 2096 19252
rect 1584 17672 1636 17678
rect 1584 17614 1636 17620
rect 2044 17264 2096 17270
rect 2044 17206 2096 17212
rect 848 17196 900 17202
rect 848 17138 900 17144
rect 860 16969 888 17138
rect 846 16960 902 16969
rect 846 16895 902 16904
rect 2056 16590 2084 17206
rect 2044 16584 2096 16590
rect 2044 16526 2096 16532
rect 1400 15496 1452 15502
rect 1400 15438 1452 15444
rect 1412 15065 1440 15438
rect 2044 15428 2096 15434
rect 2044 15370 2096 15376
rect 1398 15056 1454 15065
rect 1398 14991 1454 15000
rect 2056 14958 2084 15370
rect 2044 14952 2096 14958
rect 2044 14894 2096 14900
rect 1400 13932 1452 13938
rect 1400 13874 1452 13880
rect 1412 13705 1440 13874
rect 1398 13696 1454 13705
rect 1398 13631 1454 13640
rect 1860 12368 1912 12374
rect 1860 12310 1912 12316
rect 846 11792 902 11801
rect 846 11727 848 11736
rect 900 11727 902 11736
rect 848 11698 900 11704
rect 1872 10674 1900 12310
rect 2056 12238 2084 14894
rect 2148 12850 2176 20810
rect 2240 19854 2268 21542
rect 2424 19938 2452 22374
rect 2504 21480 2556 21486
rect 2608 21468 2636 24142
rect 3068 23798 3096 24142
rect 3056 23792 3108 23798
rect 3056 23734 3108 23740
rect 3056 23656 3108 23662
rect 3056 23598 3108 23604
rect 2780 23588 2832 23594
rect 2780 23530 2832 23536
rect 2792 21894 2820 23530
rect 3068 22642 3096 23598
rect 3160 22778 3188 27542
rect 4620 27532 4672 27538
rect 4620 27474 4672 27480
rect 3516 26988 3568 26994
rect 3516 26930 3568 26936
rect 3528 26518 3556 26930
rect 3792 26920 3844 26926
rect 3792 26862 3844 26868
rect 3884 26920 3936 26926
rect 3884 26862 3936 26868
rect 3516 26512 3568 26518
rect 3516 26454 3568 26460
rect 3804 26364 3832 26862
rect 3896 26586 3924 26862
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 3884 26580 3936 26586
rect 3884 26522 3936 26528
rect 4068 26512 4120 26518
rect 4068 26454 4120 26460
rect 3884 26376 3936 26382
rect 3804 26336 3884 26364
rect 3884 26318 3936 26324
rect 3424 25900 3476 25906
rect 3424 25842 3476 25848
rect 3436 23866 3464 25842
rect 3516 25152 3568 25158
rect 3516 25094 3568 25100
rect 3528 24274 3556 25094
rect 3608 24744 3660 24750
rect 3608 24686 3660 24692
rect 3620 24410 3648 24686
rect 3608 24404 3660 24410
rect 3608 24346 3660 24352
rect 4080 24342 4108 26454
rect 4632 26450 4660 27474
rect 5184 27470 5212 27560
rect 5448 27542 5500 27548
rect 6736 27600 6788 27606
rect 6736 27542 6788 27548
rect 5724 27532 5776 27538
rect 5724 27474 5776 27480
rect 5172 27464 5224 27470
rect 5172 27406 5224 27412
rect 5736 27402 5764 27474
rect 5908 27464 5960 27470
rect 5908 27406 5960 27412
rect 6000 27464 6052 27470
rect 6184 27464 6236 27470
rect 6052 27424 6184 27452
rect 6000 27406 6052 27412
rect 6184 27406 6236 27412
rect 5632 27396 5684 27402
rect 5632 27338 5684 27344
rect 5724 27396 5776 27402
rect 5724 27338 5776 27344
rect 5356 27328 5408 27334
rect 5356 27270 5408 27276
rect 5448 27328 5500 27334
rect 5448 27270 5500 27276
rect 5540 27328 5592 27334
rect 5540 27270 5592 27276
rect 4874 27228 5182 27237
rect 4874 27226 4880 27228
rect 4936 27226 4960 27228
rect 5016 27226 5040 27228
rect 5096 27226 5120 27228
rect 5176 27226 5182 27228
rect 4936 27174 4938 27226
rect 5118 27174 5120 27226
rect 4874 27172 4880 27174
rect 4936 27172 4960 27174
rect 5016 27172 5040 27174
rect 5096 27172 5120 27174
rect 5176 27172 5182 27174
rect 4874 27163 5182 27172
rect 5264 27124 5316 27130
rect 5264 27066 5316 27072
rect 4804 26920 4856 26926
rect 4804 26862 4856 26868
rect 4712 26784 4764 26790
rect 4712 26726 4764 26732
rect 4620 26444 4672 26450
rect 4620 26386 4672 26392
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 4620 24744 4672 24750
rect 4620 24686 4672 24692
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 4068 24336 4120 24342
rect 4068 24278 4120 24284
rect 3516 24268 3568 24274
rect 3516 24210 3568 24216
rect 4436 24132 4488 24138
rect 4632 24120 4660 24686
rect 4724 24206 4752 26726
rect 4816 26586 4844 26862
rect 4988 26784 5040 26790
rect 4988 26726 5040 26732
rect 4804 26580 4856 26586
rect 4804 26522 4856 26528
rect 5000 26382 5028 26726
rect 5172 26444 5224 26450
rect 5172 26386 5224 26392
rect 4988 26376 5040 26382
rect 4988 26318 5040 26324
rect 4804 26308 4856 26314
rect 4804 26250 4856 26256
rect 4816 24800 4844 26250
rect 5184 26246 5212 26386
rect 5276 26382 5304 27066
rect 5368 26908 5396 27270
rect 5460 27062 5488 27270
rect 5448 27056 5500 27062
rect 5448 26998 5500 27004
rect 5552 26994 5580 27270
rect 5540 26988 5592 26994
rect 5540 26930 5592 26936
rect 5448 26920 5500 26926
rect 5368 26880 5448 26908
rect 5368 26382 5396 26880
rect 5448 26862 5500 26868
rect 5552 26382 5580 26930
rect 5644 26790 5672 27338
rect 5724 26920 5776 26926
rect 5724 26862 5776 26868
rect 5632 26784 5684 26790
rect 5632 26726 5684 26732
rect 5264 26376 5316 26382
rect 5264 26318 5316 26324
rect 5356 26376 5408 26382
rect 5356 26318 5408 26324
rect 5540 26376 5592 26382
rect 5540 26318 5592 26324
rect 5172 26240 5224 26246
rect 5172 26182 5224 26188
rect 4874 26140 5182 26149
rect 4874 26138 4880 26140
rect 4936 26138 4960 26140
rect 5016 26138 5040 26140
rect 5096 26138 5120 26140
rect 5176 26138 5182 26140
rect 4936 26086 4938 26138
rect 5118 26086 5120 26138
rect 4874 26084 4880 26086
rect 4936 26084 4960 26086
rect 5016 26084 5040 26086
rect 5096 26084 5120 26086
rect 5176 26084 5182 26086
rect 4874 26075 5182 26084
rect 5736 25294 5764 26862
rect 5920 26858 5948 27406
rect 5816 26852 5868 26858
rect 5816 26794 5868 26800
rect 5908 26852 5960 26858
rect 5908 26794 5960 26800
rect 5828 26382 5856 26794
rect 6196 26790 6224 27406
rect 6748 27334 6776 27542
rect 6828 27464 6880 27470
rect 6828 27406 6880 27412
rect 6840 27334 6868 27406
rect 6736 27328 6788 27334
rect 6736 27270 6788 27276
rect 6828 27328 6880 27334
rect 6828 27270 6880 27276
rect 6644 27056 6696 27062
rect 6644 26998 6696 27004
rect 6552 26988 6604 26994
rect 6552 26930 6604 26936
rect 6184 26784 6236 26790
rect 6184 26726 6236 26732
rect 6564 26518 6592 26930
rect 6656 26518 6684 26998
rect 6932 26994 6960 27610
rect 7484 27606 7512 27950
rect 10692 27940 10744 27946
rect 10744 27900 10824 27928
rect 10692 27882 10744 27888
rect 10324 27668 10376 27674
rect 10324 27610 10376 27616
rect 7472 27600 7524 27606
rect 7472 27542 7524 27548
rect 7484 27470 7512 27542
rect 7472 27464 7524 27470
rect 7472 27406 7524 27412
rect 7656 27464 7708 27470
rect 7656 27406 7708 27412
rect 7668 27062 7696 27406
rect 10336 27334 10364 27610
rect 10508 27600 10560 27606
rect 10508 27542 10560 27548
rect 10324 27328 10376 27334
rect 10324 27270 10376 27276
rect 10416 27328 10468 27334
rect 10416 27270 10468 27276
rect 7656 27056 7708 27062
rect 10336 27033 10364 27270
rect 7656 26998 7708 27004
rect 10322 27024 10378 27033
rect 6920 26988 6972 26994
rect 6920 26930 6972 26936
rect 9128 26988 9180 26994
rect 10322 26959 10378 26968
rect 9128 26930 9180 26936
rect 6828 26920 6880 26926
rect 6828 26862 6880 26868
rect 6840 26790 6868 26862
rect 7012 26852 7064 26858
rect 7012 26794 7064 26800
rect 6828 26784 6880 26790
rect 6748 26744 6828 26772
rect 6552 26512 6604 26518
rect 6552 26454 6604 26460
rect 6644 26512 6696 26518
rect 6644 26454 6696 26460
rect 5816 26376 5868 26382
rect 5816 26318 5868 26324
rect 6644 26376 6696 26382
rect 6748 26364 6776 26744
rect 6828 26726 6880 26732
rect 6920 26784 6972 26790
rect 6920 26726 6972 26732
rect 6932 26450 6960 26726
rect 7024 26586 7052 26794
rect 7656 26784 7708 26790
rect 7656 26726 7708 26732
rect 8760 26784 8812 26790
rect 8760 26726 8812 26732
rect 7012 26580 7064 26586
rect 7012 26522 7064 26528
rect 6920 26444 6972 26450
rect 6920 26386 6972 26392
rect 7668 26382 7696 26726
rect 8772 26382 8800 26726
rect 6696 26336 6776 26364
rect 7656 26376 7708 26382
rect 6644 26318 6696 26324
rect 7656 26318 7708 26324
rect 8576 26376 8628 26382
rect 8576 26318 8628 26324
rect 8760 26376 8812 26382
rect 8760 26318 8812 26324
rect 6276 26308 6328 26314
rect 6276 26250 6328 26256
rect 5724 25288 5776 25294
rect 5724 25230 5776 25236
rect 5356 25220 5408 25226
rect 5356 25162 5408 25168
rect 4874 25052 5182 25061
rect 4874 25050 4880 25052
rect 4936 25050 4960 25052
rect 5016 25050 5040 25052
rect 5096 25050 5120 25052
rect 5176 25050 5182 25052
rect 4936 24998 4938 25050
rect 5118 24998 5120 25050
rect 4874 24996 4880 24998
rect 4936 24996 4960 24998
rect 5016 24996 5040 24998
rect 5096 24996 5120 24998
rect 5176 24996 5182 24998
rect 4874 24987 5182 24996
rect 5368 24818 5396 25162
rect 5356 24812 5408 24818
rect 4816 24772 4936 24800
rect 4804 24676 4856 24682
rect 4804 24618 4856 24624
rect 4816 24274 4844 24618
rect 4804 24268 4856 24274
rect 4804 24210 4856 24216
rect 4712 24200 4764 24206
rect 4712 24142 4764 24148
rect 4488 24092 4660 24120
rect 4436 24074 4488 24080
rect 3424 23860 3476 23866
rect 3424 23802 3476 23808
rect 3436 23594 3464 23802
rect 4448 23662 4476 24074
rect 4724 23730 4752 24142
rect 4816 23780 4844 24210
rect 4908 24138 4936 24772
rect 5356 24754 5408 24760
rect 5172 24608 5224 24614
rect 5172 24550 5224 24556
rect 5184 24206 5212 24550
rect 5368 24410 5396 24754
rect 5356 24404 5408 24410
rect 5356 24346 5408 24352
rect 5368 24256 5396 24346
rect 5368 24228 5488 24256
rect 5172 24200 5224 24206
rect 5224 24148 5396 24154
rect 5172 24142 5396 24148
rect 4896 24132 4948 24138
rect 5184 24126 5396 24142
rect 4896 24074 4948 24080
rect 5264 24064 5316 24070
rect 5264 24006 5316 24012
rect 4874 23964 5182 23973
rect 4874 23962 4880 23964
rect 4936 23962 4960 23964
rect 5016 23962 5040 23964
rect 5096 23962 5120 23964
rect 5176 23962 5182 23964
rect 4936 23910 4938 23962
rect 5118 23910 5120 23962
rect 4874 23908 4880 23910
rect 4936 23908 4960 23910
rect 5016 23908 5040 23910
rect 5096 23908 5120 23910
rect 5176 23908 5182 23910
rect 4874 23899 5182 23908
rect 4816 23752 4936 23780
rect 4620 23724 4672 23730
rect 4620 23666 4672 23672
rect 4712 23724 4764 23730
rect 4712 23666 4764 23672
rect 4436 23656 4488 23662
rect 4436 23598 4488 23604
rect 3424 23588 3476 23594
rect 3424 23530 3476 23536
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 4632 23322 4660 23666
rect 4804 23656 4856 23662
rect 4804 23598 4856 23604
rect 4620 23316 4672 23322
rect 4620 23258 4672 23264
rect 4620 23112 4672 23118
rect 4620 23054 4672 23060
rect 4712 23112 4764 23118
rect 4712 23054 4764 23060
rect 4632 22982 4660 23054
rect 4620 22976 4672 22982
rect 4620 22918 4672 22924
rect 3148 22772 3200 22778
rect 3148 22714 3200 22720
rect 3056 22636 3108 22642
rect 3056 22578 3108 22584
rect 3160 22234 3188 22714
rect 3608 22568 3660 22574
rect 3608 22510 3660 22516
rect 3240 22432 3292 22438
rect 3240 22374 3292 22380
rect 3148 22228 3200 22234
rect 3148 22170 3200 22176
rect 3252 22030 3280 22374
rect 3240 22024 3292 22030
rect 3240 21966 3292 21972
rect 3620 21962 3648 22510
rect 3884 22432 3936 22438
rect 3884 22374 3936 22380
rect 3896 22098 3924 22374
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 4160 22160 4212 22166
rect 4160 22102 4212 22108
rect 3884 22092 3936 22098
rect 3884 22034 3936 22040
rect 3700 22024 3752 22030
rect 3700 21966 3752 21972
rect 3608 21956 3660 21962
rect 3608 21898 3660 21904
rect 2780 21888 2832 21894
rect 2780 21830 2832 21836
rect 2872 21888 2924 21894
rect 2872 21830 2924 21836
rect 3424 21888 3476 21894
rect 3424 21830 3476 21836
rect 2688 21548 2740 21554
rect 2688 21490 2740 21496
rect 2556 21440 2636 21468
rect 2504 21422 2556 21428
rect 2516 20874 2544 21422
rect 2700 20942 2728 21490
rect 2688 20936 2740 20942
rect 2688 20878 2740 20884
rect 2504 20868 2556 20874
rect 2504 20810 2556 20816
rect 2700 20466 2728 20878
rect 2596 20460 2648 20466
rect 2596 20402 2648 20408
rect 2688 20460 2740 20466
rect 2688 20402 2740 20408
rect 2332 19910 2452 19938
rect 2228 19848 2280 19854
rect 2228 19790 2280 19796
rect 2240 19378 2268 19790
rect 2228 19372 2280 19378
rect 2228 19314 2280 19320
rect 2332 17882 2360 19910
rect 2412 19848 2464 19854
rect 2412 19790 2464 19796
rect 2424 19378 2452 19790
rect 2412 19372 2464 19378
rect 2412 19314 2464 19320
rect 2608 18902 2636 20402
rect 2700 19786 2728 20402
rect 2884 19854 2912 21830
rect 3436 20874 3464 21830
rect 3712 20942 3740 21966
rect 3976 21956 4028 21962
rect 3976 21898 4028 21904
rect 3988 21554 4016 21898
rect 3792 21548 3844 21554
rect 3792 21490 3844 21496
rect 3976 21548 4028 21554
rect 3976 21490 4028 21496
rect 3804 21146 3832 21490
rect 4172 21400 4200 22102
rect 4632 22094 4660 22918
rect 4724 22234 4752 23054
rect 4712 22228 4764 22234
rect 4712 22170 4764 22176
rect 4632 22066 4752 22094
rect 4724 22030 4752 22066
rect 4712 22024 4764 22030
rect 4712 21966 4764 21972
rect 4620 21888 4672 21894
rect 4620 21830 4672 21836
rect 4632 21554 4660 21830
rect 4712 21684 4764 21690
rect 4712 21626 4764 21632
rect 4620 21548 4672 21554
rect 4620 21490 4672 21496
rect 4080 21372 4200 21400
rect 3792 21140 3844 21146
rect 3792 21082 3844 21088
rect 4080 20942 4108 21372
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4632 20942 4660 21490
rect 3700 20936 3752 20942
rect 3700 20878 3752 20884
rect 4068 20936 4120 20942
rect 4620 20936 4672 20942
rect 4120 20896 4200 20924
rect 4068 20878 4120 20884
rect 3424 20868 3476 20874
rect 3424 20810 3476 20816
rect 2872 19848 2924 19854
rect 2872 19790 2924 19796
rect 2688 19780 2740 19786
rect 2688 19722 2740 19728
rect 2884 19514 2912 19790
rect 2872 19508 2924 19514
rect 2872 19450 2924 19456
rect 2688 19304 2740 19310
rect 2688 19246 2740 19252
rect 2596 18896 2648 18902
rect 2596 18838 2648 18844
rect 2608 18034 2636 18838
rect 2516 18006 2636 18034
rect 2320 17876 2372 17882
rect 2320 17818 2372 17824
rect 2516 17270 2544 18006
rect 2596 17876 2648 17882
rect 2596 17818 2648 17824
rect 2504 17264 2556 17270
rect 2504 17206 2556 17212
rect 2412 17060 2464 17066
rect 2412 17002 2464 17008
rect 2424 16794 2452 17002
rect 2412 16788 2464 16794
rect 2412 16730 2464 16736
rect 2240 16658 2360 16674
rect 2240 16652 2372 16658
rect 2240 16646 2320 16652
rect 2240 16046 2268 16646
rect 2320 16594 2372 16600
rect 2504 16584 2556 16590
rect 2608 16574 2636 17818
rect 2700 17338 2728 19246
rect 2688 17332 2740 17338
rect 2688 17274 2740 17280
rect 3240 17264 3292 17270
rect 3240 17206 3292 17212
rect 2964 16992 3016 16998
rect 2964 16934 3016 16940
rect 2976 16590 3004 16934
rect 3252 16658 3280 17206
rect 3148 16652 3200 16658
rect 3148 16594 3200 16600
rect 3240 16652 3292 16658
rect 3240 16594 3292 16600
rect 2556 16546 2636 16574
rect 2964 16584 3016 16590
rect 2504 16526 2556 16532
rect 2964 16526 3016 16532
rect 2516 16114 2544 16526
rect 2504 16108 2556 16114
rect 2504 16050 2556 16056
rect 2228 16040 2280 16046
rect 2228 15982 2280 15988
rect 2320 15904 2372 15910
rect 2320 15846 2372 15852
rect 2332 14278 2360 15846
rect 2780 15496 2832 15502
rect 2780 15438 2832 15444
rect 2792 15162 2820 15438
rect 2780 15156 2832 15162
rect 2780 15098 2832 15104
rect 3160 15026 3188 16594
rect 3252 15502 3280 16594
rect 3240 15496 3292 15502
rect 3240 15438 3292 15444
rect 3240 15360 3292 15366
rect 3240 15302 3292 15308
rect 3148 15020 3200 15026
rect 3148 14962 3200 14968
rect 3148 14816 3200 14822
rect 3148 14758 3200 14764
rect 2780 14408 2832 14414
rect 2780 14350 2832 14356
rect 2320 14272 2372 14278
rect 2320 14214 2372 14220
rect 2332 13870 2360 14214
rect 2792 14074 2820 14350
rect 2780 14068 2832 14074
rect 2780 14010 2832 14016
rect 3160 13938 3188 14758
rect 3252 14414 3280 15302
rect 3240 14408 3292 14414
rect 3240 14350 3292 14356
rect 3252 14006 3280 14350
rect 3240 14000 3292 14006
rect 3240 13942 3292 13948
rect 2688 13932 2740 13938
rect 2688 13874 2740 13880
rect 3148 13932 3200 13938
rect 3148 13874 3200 13880
rect 2320 13864 2372 13870
rect 2320 13806 2372 13812
rect 2228 13796 2280 13802
rect 2228 13738 2280 13744
rect 2240 12986 2268 13738
rect 2700 13258 2728 13874
rect 2964 13864 3016 13870
rect 2964 13806 3016 13812
rect 2976 13394 3004 13806
rect 2964 13388 3016 13394
rect 2964 13330 3016 13336
rect 3160 13326 3188 13874
rect 3148 13320 3200 13326
rect 3148 13262 3200 13268
rect 2688 13252 2740 13258
rect 2688 13194 2740 13200
rect 2228 12980 2280 12986
rect 2228 12922 2280 12928
rect 2136 12844 2188 12850
rect 2136 12786 2188 12792
rect 2412 12844 2464 12850
rect 2412 12786 2464 12792
rect 2148 12238 2176 12786
rect 2424 12306 2452 12786
rect 2700 12374 2728 13194
rect 2688 12368 2740 12374
rect 2688 12310 2740 12316
rect 2412 12300 2464 12306
rect 2412 12242 2464 12248
rect 2044 12232 2096 12238
rect 2044 12174 2096 12180
rect 2136 12232 2188 12238
rect 2136 12174 2188 12180
rect 2872 12096 2924 12102
rect 2872 12038 2924 12044
rect 1952 11688 2004 11694
rect 1952 11630 2004 11636
rect 1964 11082 1992 11630
rect 2884 11150 2912 12038
rect 2872 11144 2924 11150
rect 2872 11086 2924 11092
rect 3148 11144 3200 11150
rect 3148 11086 3200 11092
rect 1952 11076 2004 11082
rect 1952 11018 2004 11024
rect 1860 10668 1912 10674
rect 1860 10610 1912 10616
rect 1964 10606 1992 11018
rect 2884 10606 2912 11086
rect 3160 10810 3188 11086
rect 3148 10804 3200 10810
rect 3148 10746 3200 10752
rect 3436 10674 3464 20810
rect 4068 20800 4120 20806
rect 4068 20742 4120 20748
rect 4080 19938 4108 20742
rect 4172 20534 4200 20896
rect 4620 20878 4672 20884
rect 4160 20528 4212 20534
rect 4160 20470 4212 20476
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 4080 19910 4200 19938
rect 4172 19854 4200 19910
rect 4160 19848 4212 19854
rect 4160 19790 4212 19796
rect 3700 19780 3752 19786
rect 3700 19722 3752 19728
rect 3712 19310 3740 19722
rect 4724 19378 4752 21626
rect 4816 21536 4844 23598
rect 4908 22982 4936 23752
rect 5276 23186 5304 24006
rect 5368 23798 5396 24126
rect 5356 23792 5408 23798
rect 5356 23734 5408 23740
rect 5264 23180 5316 23186
rect 5264 23122 5316 23128
rect 5460 23118 5488 24228
rect 5632 23520 5684 23526
rect 5632 23462 5684 23468
rect 5540 23180 5592 23186
rect 5540 23122 5592 23128
rect 5448 23112 5500 23118
rect 5448 23054 5500 23060
rect 4896 22976 4948 22982
rect 4896 22918 4948 22924
rect 4874 22876 5182 22885
rect 4874 22874 4880 22876
rect 4936 22874 4960 22876
rect 5016 22874 5040 22876
rect 5096 22874 5120 22876
rect 5176 22874 5182 22876
rect 4936 22822 4938 22874
rect 5118 22822 5120 22874
rect 4874 22820 4880 22822
rect 4936 22820 4960 22822
rect 5016 22820 5040 22822
rect 5096 22820 5120 22822
rect 5176 22820 5182 22822
rect 4874 22811 5182 22820
rect 5552 22642 5580 23122
rect 5644 23118 5672 23462
rect 6288 23118 6316 26250
rect 6552 26240 6604 26246
rect 6552 26182 6604 26188
rect 7656 26240 7708 26246
rect 7656 26182 7708 26188
rect 6564 25362 6592 26182
rect 7668 25974 7696 26182
rect 8588 26042 8616 26318
rect 8668 26240 8720 26246
rect 8668 26182 8720 26188
rect 8576 26036 8628 26042
rect 8576 25978 8628 25984
rect 7656 25968 7708 25974
rect 7656 25910 7708 25916
rect 6552 25356 6604 25362
rect 6552 25298 6604 25304
rect 7564 25288 7616 25294
rect 7668 25276 7696 25910
rect 7932 25900 7984 25906
rect 7932 25842 7984 25848
rect 7944 25294 7972 25842
rect 8588 25294 8616 25978
rect 8680 25294 8708 26182
rect 7616 25248 7696 25276
rect 7932 25288 7984 25294
rect 7564 25230 7616 25236
rect 7932 25230 7984 25236
rect 8576 25288 8628 25294
rect 8576 25230 8628 25236
rect 8668 25288 8720 25294
rect 8668 25230 8720 25236
rect 7288 25152 7340 25158
rect 7288 25094 7340 25100
rect 7380 25152 7432 25158
rect 7380 25094 7432 25100
rect 8392 25152 8444 25158
rect 8392 25094 8444 25100
rect 7300 24206 7328 25094
rect 7392 24818 7420 25094
rect 8404 24818 8432 25094
rect 7380 24812 7432 24818
rect 7380 24754 7432 24760
rect 8116 24812 8168 24818
rect 8116 24754 8168 24760
rect 8392 24812 8444 24818
rect 8392 24754 8444 24760
rect 8128 24682 8156 24754
rect 8116 24676 8168 24682
rect 8116 24618 8168 24624
rect 8128 24410 8156 24618
rect 8576 24608 8628 24614
rect 8576 24550 8628 24556
rect 8116 24404 8168 24410
rect 8116 24346 8168 24352
rect 7472 24268 7524 24274
rect 7472 24210 7524 24216
rect 7288 24200 7340 24206
rect 7288 24142 7340 24148
rect 7300 23186 7328 24142
rect 7288 23180 7340 23186
rect 7288 23122 7340 23128
rect 7484 23118 7512 24210
rect 8588 24206 8616 24550
rect 8576 24200 8628 24206
rect 8576 24142 8628 24148
rect 8588 23798 8616 24142
rect 8576 23792 8628 23798
rect 8576 23734 8628 23740
rect 8852 23724 8904 23730
rect 8852 23666 8904 23672
rect 8864 23254 8892 23666
rect 8852 23248 8904 23254
rect 8852 23190 8904 23196
rect 8864 23118 8892 23190
rect 5632 23112 5684 23118
rect 5632 23054 5684 23060
rect 6184 23112 6236 23118
rect 6184 23054 6236 23060
rect 6276 23112 6328 23118
rect 6276 23054 6328 23060
rect 7472 23112 7524 23118
rect 7472 23054 7524 23060
rect 7932 23112 7984 23118
rect 7932 23054 7984 23060
rect 8852 23112 8904 23118
rect 8852 23054 8904 23060
rect 5540 22636 5592 22642
rect 5540 22578 5592 22584
rect 5644 22574 5672 23054
rect 6196 22642 6224 23054
rect 6184 22636 6236 22642
rect 6184 22578 6236 22584
rect 6288 22574 6316 23054
rect 7288 23044 7340 23050
rect 7288 22986 7340 22992
rect 5632 22568 5684 22574
rect 5632 22510 5684 22516
rect 6276 22568 6328 22574
rect 6276 22510 6328 22516
rect 6368 22432 6420 22438
rect 6368 22374 6420 22380
rect 4874 21788 5182 21797
rect 4874 21786 4880 21788
rect 4936 21786 4960 21788
rect 5016 21786 5040 21788
rect 5096 21786 5120 21788
rect 5176 21786 5182 21788
rect 4936 21734 4938 21786
rect 5118 21734 5120 21786
rect 4874 21732 4880 21734
rect 4936 21732 4960 21734
rect 5016 21732 5040 21734
rect 5096 21732 5120 21734
rect 5176 21732 5182 21734
rect 4874 21723 5182 21732
rect 4988 21548 5040 21554
rect 4816 21508 4988 21536
rect 4988 21490 5040 21496
rect 5000 20942 5028 21490
rect 5724 21480 5776 21486
rect 5724 21422 5776 21428
rect 5736 20942 5764 21422
rect 6380 21010 6408 22374
rect 7300 22030 7328 22986
rect 7840 22976 7892 22982
rect 7840 22918 7892 22924
rect 7852 22778 7880 22918
rect 7840 22772 7892 22778
rect 7840 22714 7892 22720
rect 7944 22438 7972 23054
rect 8024 22976 8076 22982
rect 8024 22918 8076 22924
rect 8036 22642 8064 22918
rect 8864 22710 8892 23054
rect 8852 22704 8904 22710
rect 8852 22646 8904 22652
rect 8024 22636 8076 22642
rect 8024 22578 8076 22584
rect 7380 22432 7432 22438
rect 7380 22374 7432 22380
rect 7932 22432 7984 22438
rect 7932 22374 7984 22380
rect 7392 22234 7420 22374
rect 7380 22228 7432 22234
rect 7380 22170 7432 22176
rect 7288 22024 7340 22030
rect 7288 21966 7340 21972
rect 7380 22024 7432 22030
rect 7380 21966 7432 21972
rect 7300 21486 7328 21966
rect 7392 21554 7420 21966
rect 7380 21548 7432 21554
rect 7380 21490 7432 21496
rect 7288 21480 7340 21486
rect 7288 21422 7340 21428
rect 6368 21004 6420 21010
rect 6368 20946 6420 20952
rect 4988 20936 5040 20942
rect 4988 20878 5040 20884
rect 5632 20936 5684 20942
rect 5632 20878 5684 20884
rect 5724 20936 5776 20942
rect 5724 20878 5776 20884
rect 4874 20700 5182 20709
rect 4874 20698 4880 20700
rect 4936 20698 4960 20700
rect 5016 20698 5040 20700
rect 5096 20698 5120 20700
rect 5176 20698 5182 20700
rect 4936 20646 4938 20698
rect 5118 20646 5120 20698
rect 4874 20644 4880 20646
rect 4936 20644 4960 20646
rect 5016 20644 5040 20646
rect 5096 20644 5120 20646
rect 5176 20644 5182 20646
rect 4874 20635 5182 20644
rect 4804 20460 4856 20466
rect 4804 20402 4856 20408
rect 4816 20058 4844 20402
rect 5644 20398 5672 20878
rect 5736 20466 5764 20878
rect 7104 20800 7156 20806
rect 7104 20742 7156 20748
rect 7116 20534 7144 20742
rect 7104 20528 7156 20534
rect 7104 20470 7156 20476
rect 5724 20460 5776 20466
rect 5724 20402 5776 20408
rect 5632 20392 5684 20398
rect 5632 20334 5684 20340
rect 6460 20392 6512 20398
rect 6460 20334 6512 20340
rect 4804 20052 4856 20058
rect 4804 19994 4856 20000
rect 4712 19372 4764 19378
rect 4712 19314 4764 19320
rect 3608 19304 3660 19310
rect 3608 19246 3660 19252
rect 3700 19304 3752 19310
rect 3700 19246 3752 19252
rect 3620 18902 3648 19246
rect 3608 18896 3660 18902
rect 3608 18838 3660 18844
rect 3516 18624 3568 18630
rect 3516 18566 3568 18572
rect 3528 18290 3556 18566
rect 3712 18290 3740 19246
rect 4816 19242 4844 19994
rect 5356 19848 5408 19854
rect 5356 19790 5408 19796
rect 4874 19612 5182 19621
rect 4874 19610 4880 19612
rect 4936 19610 4960 19612
rect 5016 19610 5040 19612
rect 5096 19610 5120 19612
rect 5176 19610 5182 19612
rect 4936 19558 4938 19610
rect 5118 19558 5120 19610
rect 4874 19556 4880 19558
rect 4936 19556 4960 19558
rect 5016 19556 5040 19558
rect 5096 19556 5120 19558
rect 5176 19556 5182 19558
rect 4874 19547 5182 19556
rect 5264 19304 5316 19310
rect 5264 19246 5316 19252
rect 4804 19236 4856 19242
rect 4804 19178 4856 19184
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 4816 18834 4844 19178
rect 4804 18828 4856 18834
rect 4804 18770 4856 18776
rect 5276 18766 5304 19246
rect 4436 18760 4488 18766
rect 4436 18702 4488 18708
rect 4620 18760 4672 18766
rect 4620 18702 4672 18708
rect 5264 18760 5316 18766
rect 5264 18702 5316 18708
rect 4448 18290 4476 18702
rect 4632 18290 4660 18702
rect 4874 18524 5182 18533
rect 4874 18522 4880 18524
rect 4936 18522 4960 18524
rect 5016 18522 5040 18524
rect 5096 18522 5120 18524
rect 5176 18522 5182 18524
rect 4936 18470 4938 18522
rect 5118 18470 5120 18522
rect 4874 18468 4880 18470
rect 4936 18468 4960 18470
rect 5016 18468 5040 18470
rect 5096 18468 5120 18470
rect 5176 18468 5182 18470
rect 4874 18459 5182 18468
rect 5276 18290 5304 18702
rect 3516 18284 3568 18290
rect 3516 18226 3568 18232
rect 3700 18284 3752 18290
rect 3700 18226 3752 18232
rect 4436 18284 4488 18290
rect 4436 18226 4488 18232
rect 4620 18284 4672 18290
rect 4620 18226 4672 18232
rect 5264 18284 5316 18290
rect 5264 18226 5316 18232
rect 3976 18216 4028 18222
rect 3976 18158 4028 18164
rect 3988 17202 4016 18158
rect 4632 18154 4660 18226
rect 5368 18170 5396 19790
rect 5540 19508 5592 19514
rect 5540 19450 5592 19456
rect 5552 18766 5580 19450
rect 6472 18766 6500 20334
rect 7392 19854 7420 21490
rect 8116 21480 8168 21486
rect 8116 21422 8168 21428
rect 7748 21004 7800 21010
rect 7748 20946 7800 20952
rect 7564 20460 7616 20466
rect 7564 20402 7616 20408
rect 7576 19854 7604 20402
rect 7760 20398 7788 20946
rect 7748 20392 7800 20398
rect 7748 20334 7800 20340
rect 7760 19922 7788 20334
rect 7748 19916 7800 19922
rect 7748 19858 7800 19864
rect 8128 19854 8156 21422
rect 8392 20596 8444 20602
rect 8392 20538 8444 20544
rect 7380 19848 7432 19854
rect 7380 19790 7432 19796
rect 7564 19848 7616 19854
rect 7564 19790 7616 19796
rect 8116 19848 8168 19854
rect 8116 19790 8168 19796
rect 7576 19242 7604 19790
rect 7840 19712 7892 19718
rect 7840 19654 7892 19660
rect 7852 19378 7880 19654
rect 8128 19378 8156 19790
rect 8404 19786 8432 20538
rect 9140 19990 9168 26930
rect 9864 26920 9916 26926
rect 9864 26862 9916 26868
rect 9772 26784 9824 26790
rect 9772 26726 9824 26732
rect 9784 26382 9812 26726
rect 9876 26586 9904 26862
rect 10428 26858 10456 27270
rect 9956 26852 10008 26858
rect 9956 26794 10008 26800
rect 10416 26852 10468 26858
rect 10416 26794 10468 26800
rect 9968 26586 9996 26794
rect 10232 26784 10284 26790
rect 10232 26726 10284 26732
rect 9864 26580 9916 26586
rect 9864 26522 9916 26528
rect 9956 26580 10008 26586
rect 9956 26522 10008 26528
rect 10244 26518 10272 26726
rect 10232 26512 10284 26518
rect 10232 26454 10284 26460
rect 10520 26382 10548 27542
rect 10796 27470 10824 27900
rect 11072 27674 11100 28018
rect 11152 27940 11204 27946
rect 11152 27882 11204 27888
rect 11060 27668 11112 27674
rect 11060 27610 11112 27616
rect 10968 27600 11020 27606
rect 10968 27542 11020 27548
rect 10600 27464 10652 27470
rect 10600 27406 10652 27412
rect 10784 27464 10836 27470
rect 10784 27406 10836 27412
rect 10612 27334 10640 27406
rect 10600 27328 10652 27334
rect 10600 27270 10652 27276
rect 10612 26994 10640 27270
rect 10796 26994 10824 27406
rect 10980 26994 11008 27542
rect 11072 27130 11100 27610
rect 11060 27124 11112 27130
rect 11060 27066 11112 27072
rect 11058 27024 11114 27033
rect 10600 26988 10652 26994
rect 10600 26930 10652 26936
rect 10784 26988 10836 26994
rect 10784 26930 10836 26936
rect 10968 26988 11020 26994
rect 11058 26959 11060 26968
rect 10968 26930 11020 26936
rect 11112 26959 11114 26968
rect 11060 26930 11112 26936
rect 10600 26784 10652 26790
rect 10600 26726 10652 26732
rect 10612 26602 10640 26726
rect 10612 26574 10732 26602
rect 11164 26586 11192 27882
rect 11244 27872 11296 27878
rect 11244 27814 11296 27820
rect 11256 27470 11284 27814
rect 11716 27470 11744 28018
rect 15856 28014 15884 28494
rect 15844 28008 15896 28014
rect 15844 27950 15896 27956
rect 16960 27606 16988 28494
rect 17144 28218 17172 28494
rect 17408 28484 17460 28490
rect 17408 28426 17460 28432
rect 17224 28416 17276 28422
rect 17224 28358 17276 28364
rect 17132 28212 17184 28218
rect 17132 28154 17184 28160
rect 17236 27606 17264 28358
rect 16948 27600 17000 27606
rect 16948 27542 17000 27548
rect 17224 27600 17276 27606
rect 17224 27542 17276 27548
rect 11244 27464 11296 27470
rect 11244 27406 11296 27412
rect 11704 27464 11756 27470
rect 11704 27406 11756 27412
rect 11888 27464 11940 27470
rect 11888 27406 11940 27412
rect 16948 27464 17000 27470
rect 16948 27406 17000 27412
rect 11256 26790 11284 27406
rect 11716 26790 11744 27406
rect 11244 26784 11296 26790
rect 11244 26726 11296 26732
rect 11520 26784 11572 26790
rect 11520 26726 11572 26732
rect 11704 26784 11756 26790
rect 11704 26726 11756 26732
rect 10704 26382 10732 26574
rect 11152 26580 11204 26586
rect 11152 26522 11204 26528
rect 11532 26382 11560 26726
rect 11716 26518 11744 26726
rect 11704 26512 11756 26518
rect 11704 26454 11756 26460
rect 11900 26450 11928 27406
rect 11980 27328 12032 27334
rect 11980 27270 12032 27276
rect 11992 27062 12020 27270
rect 12348 27124 12400 27130
rect 12348 27066 12400 27072
rect 11980 27056 12032 27062
rect 11980 26998 12032 27004
rect 12256 26580 12308 26586
rect 12256 26522 12308 26528
rect 11888 26444 11940 26450
rect 11888 26386 11940 26392
rect 12268 26382 12296 26522
rect 9772 26376 9824 26382
rect 9772 26318 9824 26324
rect 10232 26376 10284 26382
rect 10508 26376 10560 26382
rect 10284 26336 10508 26364
rect 10232 26318 10284 26324
rect 10508 26318 10560 26324
rect 10692 26376 10744 26382
rect 10692 26318 10744 26324
rect 11520 26376 11572 26382
rect 11520 26318 11572 26324
rect 12164 26376 12216 26382
rect 12164 26318 12216 26324
rect 12256 26376 12308 26382
rect 12256 26318 12308 26324
rect 10520 26246 10548 26318
rect 12072 26308 12124 26314
rect 12072 26250 12124 26256
rect 9404 26240 9456 26246
rect 9404 26182 9456 26188
rect 10048 26240 10100 26246
rect 10048 26182 10100 26188
rect 10416 26240 10468 26246
rect 10416 26182 10468 26188
rect 10508 26240 10560 26246
rect 10508 26182 10560 26188
rect 9416 25294 9444 26182
rect 10060 25974 10088 26182
rect 10048 25968 10100 25974
rect 10048 25910 10100 25916
rect 10324 25968 10376 25974
rect 10324 25910 10376 25916
rect 10048 25424 10100 25430
rect 10048 25366 10100 25372
rect 9404 25288 9456 25294
rect 9404 25230 9456 25236
rect 9496 25152 9548 25158
rect 9496 25094 9548 25100
rect 9508 24818 9536 25094
rect 10060 24886 10088 25366
rect 10048 24880 10100 24886
rect 10048 24822 10100 24828
rect 10336 24818 10364 25910
rect 10428 25906 10456 26182
rect 10416 25900 10468 25906
rect 10416 25842 10468 25848
rect 10428 25294 10456 25842
rect 10508 25696 10560 25702
rect 10508 25638 10560 25644
rect 10520 25430 10548 25638
rect 10508 25424 10560 25430
rect 10508 25366 10560 25372
rect 10416 25288 10468 25294
rect 10416 25230 10468 25236
rect 11980 25288 12032 25294
rect 11980 25230 12032 25236
rect 10508 25152 10560 25158
rect 10508 25094 10560 25100
rect 10520 24818 10548 25094
rect 11992 24954 12020 25230
rect 11980 24948 12032 24954
rect 11980 24890 12032 24896
rect 12084 24818 12112 26250
rect 12176 24954 12204 26318
rect 12360 26246 12388 27066
rect 16960 27062 16988 27406
rect 17420 27130 17448 28426
rect 17776 28416 17828 28422
rect 17776 28358 17828 28364
rect 17788 27606 17816 28358
rect 17776 27600 17828 27606
rect 17776 27542 17828 27548
rect 17408 27124 17460 27130
rect 17408 27066 17460 27072
rect 12992 27056 13044 27062
rect 12992 26998 13044 27004
rect 16948 27056 17000 27062
rect 16948 26998 17000 27004
rect 12716 26988 12768 26994
rect 12716 26930 12768 26936
rect 12532 26784 12584 26790
rect 12532 26726 12584 26732
rect 12544 26586 12572 26726
rect 12532 26580 12584 26586
rect 12452 26540 12532 26568
rect 12348 26240 12400 26246
rect 12348 26182 12400 26188
rect 12452 25294 12480 26540
rect 12532 26522 12584 26528
rect 12728 26382 12756 26930
rect 12716 26376 12768 26382
rect 12716 26318 12768 26324
rect 12808 26376 12860 26382
rect 12808 26318 12860 26324
rect 12532 26240 12584 26246
rect 12532 26182 12584 26188
rect 12544 25906 12572 26182
rect 12728 26042 12756 26318
rect 12716 26036 12768 26042
rect 12716 25978 12768 25984
rect 12532 25900 12584 25906
rect 12532 25842 12584 25848
rect 12716 25900 12768 25906
rect 12716 25842 12768 25848
rect 12728 25294 12756 25842
rect 12348 25288 12400 25294
rect 12348 25230 12400 25236
rect 12440 25288 12492 25294
rect 12440 25230 12492 25236
rect 12716 25288 12768 25294
rect 12716 25230 12768 25236
rect 12164 24948 12216 24954
rect 12164 24890 12216 24896
rect 9496 24812 9548 24818
rect 9496 24754 9548 24760
rect 10324 24812 10376 24818
rect 10324 24754 10376 24760
rect 10508 24812 10560 24818
rect 10508 24754 10560 24760
rect 11796 24812 11848 24818
rect 11796 24754 11848 24760
rect 12072 24812 12124 24818
rect 12072 24754 12124 24760
rect 9404 24608 9456 24614
rect 9404 24550 9456 24556
rect 9312 24336 9364 24342
rect 9312 24278 9364 24284
rect 9324 23254 9352 24278
rect 9416 24206 9444 24550
rect 9508 24206 9536 24754
rect 10416 24744 10468 24750
rect 10416 24686 10468 24692
rect 9956 24608 10008 24614
rect 9956 24550 10008 24556
rect 10324 24608 10376 24614
rect 10324 24550 10376 24556
rect 9404 24200 9456 24206
rect 9404 24142 9456 24148
rect 9496 24200 9548 24206
rect 9496 24142 9548 24148
rect 9772 24200 9824 24206
rect 9772 24142 9824 24148
rect 9864 24200 9916 24206
rect 9864 24142 9916 24148
rect 9416 23730 9444 24142
rect 9784 23798 9812 24142
rect 9772 23792 9824 23798
rect 9772 23734 9824 23740
rect 9404 23724 9456 23730
rect 9404 23666 9456 23672
rect 9312 23248 9364 23254
rect 9312 23190 9364 23196
rect 9324 23118 9352 23190
rect 9312 23112 9364 23118
rect 9496 23112 9548 23118
rect 9312 23054 9364 23060
rect 9416 23072 9496 23100
rect 9220 22636 9272 22642
rect 9220 22578 9272 22584
rect 9232 22030 9260 22578
rect 9324 22438 9352 23054
rect 9416 22710 9444 23072
rect 9496 23054 9548 23060
rect 9772 22976 9824 22982
rect 9772 22918 9824 22924
rect 9404 22704 9456 22710
rect 9404 22646 9456 22652
rect 9312 22432 9364 22438
rect 9312 22374 9364 22380
rect 9416 22030 9444 22646
rect 9784 22642 9812 22918
rect 9876 22710 9904 24142
rect 9968 23118 9996 24550
rect 10336 23594 10364 24550
rect 10428 24206 10456 24686
rect 10416 24200 10468 24206
rect 10416 24142 10468 24148
rect 10428 23866 10456 24142
rect 11808 24138 11836 24754
rect 11980 24744 12032 24750
rect 11980 24686 12032 24692
rect 11992 24410 12020 24686
rect 11980 24404 12032 24410
rect 11980 24346 12032 24352
rect 12084 24138 12112 24754
rect 11796 24132 11848 24138
rect 11796 24074 11848 24080
rect 12072 24132 12124 24138
rect 12072 24074 12124 24080
rect 10416 23860 10468 23866
rect 10416 23802 10468 23808
rect 10324 23588 10376 23594
rect 10324 23530 10376 23536
rect 11808 23322 11836 24074
rect 12176 23662 12204 24890
rect 12360 24682 12388 25230
rect 12348 24676 12400 24682
rect 12348 24618 12400 24624
rect 12360 24206 12388 24618
rect 12440 24608 12492 24614
rect 12440 24550 12492 24556
rect 12348 24200 12400 24206
rect 12348 24142 12400 24148
rect 12256 23724 12308 23730
rect 12360 23712 12388 24142
rect 12452 23866 12480 24550
rect 12716 24200 12768 24206
rect 12820 24188 12848 26318
rect 13004 26246 13032 26998
rect 17880 26858 17908 28494
rect 17972 27334 18000 28562
rect 18052 27940 18104 27946
rect 18052 27882 18104 27888
rect 17960 27328 18012 27334
rect 17960 27270 18012 27276
rect 18064 27130 18092 27882
rect 18156 27130 18184 28630
rect 19984 28620 20036 28626
rect 19984 28562 20036 28568
rect 19064 28552 19116 28558
rect 19064 28494 19116 28500
rect 19432 28552 19484 28558
rect 19432 28494 19484 28500
rect 19892 28552 19944 28558
rect 19892 28494 19944 28500
rect 18696 28416 18748 28422
rect 18696 28358 18748 28364
rect 18708 28082 18736 28358
rect 19076 28218 19104 28494
rect 19064 28212 19116 28218
rect 19064 28154 19116 28160
rect 18604 28076 18656 28082
rect 18604 28018 18656 28024
rect 18696 28076 18748 28082
rect 18696 28018 18748 28024
rect 18236 27668 18288 27674
rect 18236 27610 18288 27616
rect 18248 27334 18276 27610
rect 18616 27606 18644 28018
rect 18604 27600 18656 27606
rect 18604 27542 18656 27548
rect 18708 27538 18736 28018
rect 19064 28008 19116 28014
rect 19064 27950 19116 27956
rect 18788 27872 18840 27878
rect 18788 27814 18840 27820
rect 18800 27674 18828 27814
rect 18788 27668 18840 27674
rect 18788 27610 18840 27616
rect 18696 27532 18748 27538
rect 18696 27474 18748 27480
rect 18788 27532 18840 27538
rect 18788 27474 18840 27480
rect 18512 27464 18564 27470
rect 18512 27406 18564 27412
rect 18236 27328 18288 27334
rect 18236 27270 18288 27276
rect 18328 27328 18380 27334
rect 18328 27270 18380 27276
rect 18052 27124 18104 27130
rect 18052 27066 18104 27072
rect 18144 27124 18196 27130
rect 18144 27066 18196 27072
rect 17960 26988 18012 26994
rect 17960 26930 18012 26936
rect 17972 26858 18000 26930
rect 17868 26852 17920 26858
rect 17868 26794 17920 26800
rect 17960 26852 18012 26858
rect 17960 26794 18012 26800
rect 18340 26790 18368 27270
rect 18524 27062 18552 27406
rect 18512 27056 18564 27062
rect 18512 26998 18564 27004
rect 18524 26790 18552 26998
rect 18708 26994 18736 27474
rect 18696 26988 18748 26994
rect 18696 26930 18748 26936
rect 18800 26858 18828 27474
rect 19076 27334 19104 27950
rect 19156 27940 19208 27946
rect 19156 27882 19208 27888
rect 19168 27402 19196 27882
rect 19248 27668 19300 27674
rect 19248 27610 19300 27616
rect 19260 27470 19288 27610
rect 19248 27464 19300 27470
rect 19248 27406 19300 27412
rect 19156 27396 19208 27402
rect 19156 27338 19208 27344
rect 19064 27328 19116 27334
rect 19064 27270 19116 27276
rect 19260 26858 19288 27406
rect 19444 27130 19472 28494
rect 19524 28076 19576 28082
rect 19524 28018 19576 28024
rect 19536 27334 19564 28018
rect 19616 28008 19668 28014
rect 19616 27950 19668 27956
rect 19628 27470 19656 27950
rect 19708 27940 19760 27946
rect 19760 27900 19840 27928
rect 19708 27882 19760 27888
rect 19616 27464 19668 27470
rect 19616 27406 19668 27412
rect 19524 27328 19576 27334
rect 19524 27270 19576 27276
rect 19432 27124 19484 27130
rect 19432 27066 19484 27072
rect 19536 26994 19564 27270
rect 19524 26988 19576 26994
rect 19524 26930 19576 26936
rect 18788 26852 18840 26858
rect 18788 26794 18840 26800
rect 19248 26852 19300 26858
rect 19248 26794 19300 26800
rect 18328 26784 18380 26790
rect 18328 26726 18380 26732
rect 18512 26784 18564 26790
rect 18512 26726 18564 26732
rect 18340 26586 18368 26726
rect 18328 26580 18380 26586
rect 18328 26522 18380 26528
rect 19628 26450 19656 27406
rect 19812 27402 19840 27900
rect 19904 27674 19932 28494
rect 19996 28014 20024 28562
rect 20444 28552 20496 28558
rect 20444 28494 20496 28500
rect 21364 28552 21416 28558
rect 21364 28494 21416 28500
rect 22284 28552 22336 28558
rect 22284 28494 22336 28500
rect 22652 28552 22704 28558
rect 22652 28494 22704 28500
rect 23296 28552 23348 28558
rect 23296 28494 23348 28500
rect 23940 28552 23992 28558
rect 23940 28494 23992 28500
rect 24584 28552 24636 28558
rect 24584 28494 24636 28500
rect 24952 28552 25004 28558
rect 24952 28494 25004 28500
rect 25872 28552 25924 28558
rect 25872 28494 25924 28500
rect 26056 28552 26108 28558
rect 26056 28494 26108 28500
rect 26792 28552 26844 28558
rect 26792 28494 26844 28500
rect 20076 28416 20128 28422
rect 20076 28358 20128 28364
rect 20088 28082 20116 28358
rect 20456 28218 20484 28494
rect 20444 28212 20496 28218
rect 20444 28154 20496 28160
rect 20076 28076 20128 28082
rect 20076 28018 20128 28024
rect 20352 28076 20404 28082
rect 20352 28018 20404 28024
rect 19984 28008 20036 28014
rect 19984 27950 20036 27956
rect 19892 27668 19944 27674
rect 19996 27656 20024 27950
rect 20076 27668 20128 27674
rect 19996 27628 20076 27656
rect 19892 27610 19944 27616
rect 20076 27610 20128 27616
rect 19800 27396 19852 27402
rect 19800 27338 19852 27344
rect 19812 26994 19840 27338
rect 19984 27056 20036 27062
rect 19982 27024 19984 27033
rect 20036 27024 20038 27033
rect 19800 26988 19852 26994
rect 19982 26959 20038 26968
rect 19800 26930 19852 26936
rect 19996 26926 20024 26959
rect 19984 26920 20036 26926
rect 19984 26862 20036 26868
rect 19616 26444 19668 26450
rect 19616 26386 19668 26392
rect 19996 26382 20024 26862
rect 13084 26376 13136 26382
rect 13084 26318 13136 26324
rect 19984 26376 20036 26382
rect 19984 26318 20036 26324
rect 12992 26240 13044 26246
rect 12992 26182 13044 26188
rect 12900 25152 12952 25158
rect 12900 25094 12952 25100
rect 12768 24160 12848 24188
rect 12716 24142 12768 24148
rect 12440 23860 12492 23866
rect 12492 23820 12572 23848
rect 12440 23802 12492 23808
rect 12440 23724 12492 23730
rect 12360 23684 12440 23712
rect 12256 23666 12308 23672
rect 12440 23666 12492 23672
rect 12164 23656 12216 23662
rect 12164 23598 12216 23604
rect 12164 23520 12216 23526
rect 12164 23462 12216 23468
rect 11796 23316 11848 23322
rect 11796 23258 11848 23264
rect 10324 23180 10376 23186
rect 10324 23122 10376 23128
rect 9956 23112 10008 23118
rect 9956 23054 10008 23060
rect 10232 23112 10284 23118
rect 10232 23054 10284 23060
rect 10244 22778 10272 23054
rect 10232 22772 10284 22778
rect 10232 22714 10284 22720
rect 9864 22704 9916 22710
rect 9864 22646 9916 22652
rect 10336 22642 10364 23122
rect 10508 23112 10560 23118
rect 10508 23054 10560 23060
rect 10520 22710 10548 23054
rect 10508 22704 10560 22710
rect 10508 22646 10560 22652
rect 9772 22636 9824 22642
rect 9772 22578 9824 22584
rect 10048 22636 10100 22642
rect 10048 22578 10100 22584
rect 10324 22636 10376 22642
rect 10324 22578 10376 22584
rect 9784 22030 9812 22578
rect 10060 22438 10088 22578
rect 10048 22432 10100 22438
rect 10048 22374 10100 22380
rect 9220 22024 9272 22030
rect 9220 21966 9272 21972
rect 9404 22024 9456 22030
rect 9404 21966 9456 21972
rect 9772 22024 9824 22030
rect 9772 21966 9824 21972
rect 9128 19984 9180 19990
rect 9128 19926 9180 19932
rect 8392 19780 8444 19786
rect 8392 19722 8444 19728
rect 8404 19378 8432 19722
rect 7840 19372 7892 19378
rect 7840 19314 7892 19320
rect 8116 19372 8168 19378
rect 8392 19372 8444 19378
rect 8168 19332 8340 19360
rect 8116 19314 8168 19320
rect 7564 19236 7616 19242
rect 7564 19178 7616 19184
rect 5540 18760 5592 18766
rect 5540 18702 5592 18708
rect 6460 18760 6512 18766
rect 6460 18702 6512 18708
rect 6472 18358 6500 18702
rect 6552 18692 6604 18698
rect 6552 18634 6604 18640
rect 6460 18352 6512 18358
rect 6460 18294 6512 18300
rect 6564 18290 6592 18634
rect 7576 18290 7604 19178
rect 7932 19168 7984 19174
rect 7932 19110 7984 19116
rect 8208 19168 8260 19174
rect 8208 19110 8260 19116
rect 7944 18834 7972 19110
rect 7932 18828 7984 18834
rect 7932 18770 7984 18776
rect 7748 18692 7800 18698
rect 7748 18634 7800 18640
rect 6552 18284 6604 18290
rect 6552 18226 6604 18232
rect 7380 18284 7432 18290
rect 7380 18226 7432 18232
rect 7564 18284 7616 18290
rect 7564 18226 7616 18232
rect 4620 18148 4672 18154
rect 4620 18090 4672 18096
rect 5276 18142 5396 18170
rect 5816 18216 5868 18222
rect 5816 18158 5868 18164
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 3792 17196 3844 17202
rect 3792 17138 3844 17144
rect 3976 17196 4028 17202
rect 3976 17138 4028 17144
rect 3804 16658 3832 17138
rect 3884 16992 3936 16998
rect 3884 16934 3936 16940
rect 3792 16652 3844 16658
rect 3792 16594 3844 16600
rect 3896 16114 3924 16934
rect 3988 16590 4016 17138
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4632 16726 4660 18090
rect 4874 17436 5182 17445
rect 4874 17434 4880 17436
rect 4936 17434 4960 17436
rect 5016 17434 5040 17436
rect 5096 17434 5120 17436
rect 5176 17434 5182 17436
rect 4936 17382 4938 17434
rect 5118 17382 5120 17434
rect 4874 17380 4880 17382
rect 4936 17380 4960 17382
rect 5016 17380 5040 17382
rect 5096 17380 5120 17382
rect 5176 17380 5182 17382
rect 4874 17371 5182 17380
rect 4620 16720 4672 16726
rect 4620 16662 4672 16668
rect 3976 16584 4028 16590
rect 3976 16526 4028 16532
rect 4528 16584 4580 16590
rect 4528 16526 4580 16532
rect 3884 16108 3936 16114
rect 3884 16050 3936 16056
rect 4540 16046 4568 16526
rect 4620 16448 4672 16454
rect 4620 16390 4672 16396
rect 4632 16114 4660 16390
rect 4874 16348 5182 16357
rect 4874 16346 4880 16348
rect 4936 16346 4960 16348
rect 5016 16346 5040 16348
rect 5096 16346 5120 16348
rect 5176 16346 5182 16348
rect 4936 16294 4938 16346
rect 5118 16294 5120 16346
rect 4874 16292 4880 16294
rect 4936 16292 4960 16294
rect 5016 16292 5040 16294
rect 5096 16292 5120 16294
rect 5176 16292 5182 16294
rect 4874 16283 5182 16292
rect 4620 16108 4672 16114
rect 4620 16050 4672 16056
rect 4896 16108 4948 16114
rect 4896 16050 4948 16056
rect 4528 16040 4580 16046
rect 4528 15982 4580 15988
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4632 15570 4660 16050
rect 4620 15564 4672 15570
rect 4620 15506 4672 15512
rect 4908 15502 4936 16050
rect 4896 15496 4948 15502
rect 4632 15444 4896 15450
rect 4632 15438 4948 15444
rect 4632 15422 4936 15438
rect 4632 14822 4660 15422
rect 4804 15360 4856 15366
rect 4804 15302 4856 15308
rect 4816 14890 4844 15302
rect 4874 15260 5182 15269
rect 4874 15258 4880 15260
rect 4936 15258 4960 15260
rect 5016 15258 5040 15260
rect 5096 15258 5120 15260
rect 5176 15258 5182 15260
rect 4936 15206 4938 15258
rect 5118 15206 5120 15258
rect 4874 15204 4880 15206
rect 4936 15204 4960 15206
rect 5016 15204 5040 15206
rect 5096 15204 5120 15206
rect 5176 15204 5182 15206
rect 4874 15195 5182 15204
rect 4804 14884 4856 14890
rect 4804 14826 4856 14832
rect 4620 14816 4672 14822
rect 4620 14758 4672 14764
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4252 14476 4304 14482
rect 4252 14418 4304 14424
rect 3608 14408 3660 14414
rect 3608 14350 3660 14356
rect 4160 14408 4212 14414
rect 4160 14350 4212 14356
rect 3620 14074 3648 14350
rect 3700 14272 3752 14278
rect 3700 14214 3752 14220
rect 3608 14068 3660 14074
rect 3608 14010 3660 14016
rect 3712 13938 3740 14214
rect 4172 13938 4200 14350
rect 4264 13938 4292 14418
rect 4632 14414 4660 14758
rect 4712 14544 4764 14550
rect 4712 14486 4764 14492
rect 4620 14408 4672 14414
rect 4620 14350 4672 14356
rect 3700 13932 3752 13938
rect 3700 13874 3752 13880
rect 4160 13932 4212 13938
rect 4160 13874 4212 13880
rect 4252 13932 4304 13938
rect 4252 13874 4304 13880
rect 4620 13728 4672 13734
rect 4620 13670 4672 13676
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4632 13326 4660 13670
rect 4724 13394 4752 14486
rect 4816 14414 4844 14826
rect 4804 14408 4856 14414
rect 4804 14350 4856 14356
rect 4874 14172 5182 14181
rect 4874 14170 4880 14172
rect 4936 14170 4960 14172
rect 5016 14170 5040 14172
rect 5096 14170 5120 14172
rect 5176 14170 5182 14172
rect 4936 14118 4938 14170
rect 5118 14118 5120 14170
rect 4874 14116 4880 14118
rect 4936 14116 4960 14118
rect 5016 14116 5040 14118
rect 5096 14116 5120 14118
rect 5176 14116 5182 14118
rect 4874 14107 5182 14116
rect 5276 14090 5304 18142
rect 5632 17128 5684 17134
rect 5632 17070 5684 17076
rect 5356 16720 5408 16726
rect 5356 16662 5408 16668
rect 5368 16114 5396 16662
rect 5644 16454 5672 17070
rect 5828 16590 5856 18158
rect 7392 17678 7420 18226
rect 7760 18222 7788 18634
rect 7944 18426 7972 18770
rect 8220 18766 8248 19110
rect 8312 18766 8340 19332
rect 8392 19314 8444 19320
rect 8944 19372 8996 19378
rect 8944 19314 8996 19320
rect 8208 18760 8260 18766
rect 8208 18702 8260 18708
rect 8300 18760 8352 18766
rect 8300 18702 8352 18708
rect 8404 18698 8432 19314
rect 8956 18766 8984 19314
rect 8944 18760 8996 18766
rect 8944 18702 8996 18708
rect 8392 18692 8444 18698
rect 8392 18634 8444 18640
rect 8300 18624 8352 18630
rect 8300 18566 8352 18572
rect 7932 18420 7984 18426
rect 7932 18362 7984 18368
rect 7748 18216 7800 18222
rect 7748 18158 7800 18164
rect 7840 18216 7892 18222
rect 7840 18158 7892 18164
rect 7760 17678 7788 18158
rect 7380 17672 7432 17678
rect 7380 17614 7432 17620
rect 7656 17672 7708 17678
rect 7656 17614 7708 17620
rect 7748 17672 7800 17678
rect 7748 17614 7800 17620
rect 7288 17196 7340 17202
rect 7288 17138 7340 17144
rect 6920 17128 6972 17134
rect 6920 17070 6972 17076
rect 5816 16584 5868 16590
rect 5816 16526 5868 16532
rect 6932 16522 6960 17070
rect 6920 16516 6972 16522
rect 6920 16458 6972 16464
rect 5632 16448 5684 16454
rect 5632 16390 5684 16396
rect 6932 16250 6960 16458
rect 6920 16244 6972 16250
rect 6920 16186 6972 16192
rect 7300 16114 7328 17138
rect 7564 16516 7616 16522
rect 7564 16458 7616 16464
rect 5356 16108 5408 16114
rect 5356 16050 5408 16056
rect 7288 16108 7340 16114
rect 7288 16050 7340 16056
rect 5368 15502 5396 16050
rect 7576 15706 7604 16458
rect 7564 15700 7616 15706
rect 7564 15642 7616 15648
rect 5356 15496 5408 15502
rect 5356 15438 5408 15444
rect 5368 15094 5396 15438
rect 5356 15088 5408 15094
rect 5356 15030 5408 15036
rect 5368 14260 5396 15030
rect 7668 15026 7696 17614
rect 7852 16794 7880 18158
rect 8312 17814 8340 18566
rect 8668 18148 8720 18154
rect 8668 18090 8720 18096
rect 8300 17808 8352 17814
rect 8300 17750 8352 17756
rect 8576 17604 8628 17610
rect 8576 17546 8628 17552
rect 8588 17202 8616 17546
rect 8024 17196 8076 17202
rect 8024 17138 8076 17144
rect 8576 17196 8628 17202
rect 8576 17138 8628 17144
rect 8036 17066 8064 17138
rect 8024 17060 8076 17066
rect 8024 17002 8076 17008
rect 7840 16788 7892 16794
rect 7840 16730 7892 16736
rect 8036 16590 8064 17002
rect 8024 16584 8076 16590
rect 7944 16544 8024 16572
rect 7944 15502 7972 16544
rect 8484 16584 8536 16590
rect 8024 16526 8076 16532
rect 8404 16544 8484 16572
rect 8300 16516 8352 16522
rect 8300 16458 8352 16464
rect 8208 16108 8260 16114
rect 8208 16050 8260 16056
rect 7932 15496 7984 15502
rect 7932 15438 7984 15444
rect 7656 15020 7708 15026
rect 7656 14962 7708 14968
rect 5448 14952 5500 14958
rect 5448 14894 5500 14900
rect 5460 14414 5488 14894
rect 6184 14816 6236 14822
rect 6184 14758 6236 14764
rect 5908 14476 5960 14482
rect 5908 14418 5960 14424
rect 5448 14408 5500 14414
rect 5448 14350 5500 14356
rect 5368 14232 5488 14260
rect 5276 14062 5396 14090
rect 4804 13932 4856 13938
rect 4804 13874 4856 13880
rect 4712 13388 4764 13394
rect 4712 13330 4764 13336
rect 4620 13320 4672 13326
rect 4620 13262 4672 13268
rect 3792 13184 3844 13190
rect 3792 13126 3844 13132
rect 3804 11694 3832 13126
rect 4712 12844 4764 12850
rect 4712 12786 4764 12792
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4528 11892 4580 11898
rect 4528 11834 4580 11840
rect 4540 11762 4568 11834
rect 4724 11830 4752 12786
rect 4816 11830 4844 13874
rect 5264 13184 5316 13190
rect 5264 13126 5316 13132
rect 4874 13084 5182 13093
rect 4874 13082 4880 13084
rect 4936 13082 4960 13084
rect 5016 13082 5040 13084
rect 5096 13082 5120 13084
rect 5176 13082 5182 13084
rect 4936 13030 4938 13082
rect 5118 13030 5120 13082
rect 4874 13028 4880 13030
rect 4936 13028 4960 13030
rect 5016 13028 5040 13030
rect 5096 13028 5120 13030
rect 5176 13028 5182 13030
rect 4874 13019 5182 13028
rect 5276 12986 5304 13126
rect 5264 12980 5316 12986
rect 5264 12922 5316 12928
rect 5368 12434 5396 14062
rect 5276 12406 5396 12434
rect 4874 11996 5182 12005
rect 4874 11994 4880 11996
rect 4936 11994 4960 11996
rect 5016 11994 5040 11996
rect 5096 11994 5120 11996
rect 5176 11994 5182 11996
rect 4936 11942 4938 11994
rect 5118 11942 5120 11994
rect 4874 11940 4880 11942
rect 4936 11940 4960 11942
rect 5016 11940 5040 11942
rect 5096 11940 5120 11942
rect 5176 11940 5182 11942
rect 4874 11931 5182 11940
rect 4712 11824 4764 11830
rect 4712 11766 4764 11772
rect 4804 11824 4856 11830
rect 4804 11766 4856 11772
rect 4528 11756 4580 11762
rect 4580 11716 4660 11744
rect 4528 11698 4580 11704
rect 3792 11688 3844 11694
rect 3792 11630 3844 11636
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4632 11354 4660 11716
rect 4620 11348 4672 11354
rect 4620 11290 4672 11296
rect 4816 11218 4844 11766
rect 4896 11756 4948 11762
rect 4896 11698 4948 11704
rect 4908 11218 4936 11698
rect 4804 11212 4856 11218
rect 4804 11154 4856 11160
rect 4896 11212 4948 11218
rect 4896 11154 4948 11160
rect 4160 11144 4212 11150
rect 4160 11086 4212 11092
rect 3424 10668 3476 10674
rect 3424 10610 3476 10616
rect 1952 10600 2004 10606
rect 1952 10542 2004 10548
rect 2872 10600 2924 10606
rect 2872 10542 2924 10548
rect 2688 10532 2740 10538
rect 2688 10474 2740 10480
rect 2700 10130 2728 10474
rect 2688 10124 2740 10130
rect 2688 10066 2740 10072
rect 3436 10062 3464 10610
rect 4068 10464 4120 10470
rect 4172 10452 4200 11086
rect 4712 11008 4764 11014
rect 4712 10950 4764 10956
rect 4120 10424 4200 10452
rect 4068 10406 4120 10412
rect 4080 10130 4108 10406
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4620 10192 4672 10198
rect 4620 10134 4672 10140
rect 4068 10124 4120 10130
rect 4068 10066 4120 10072
rect 3424 10056 3476 10062
rect 3424 9998 3476 10004
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4632 7954 4660 10134
rect 4724 10062 4752 10950
rect 4874 10908 5182 10917
rect 4874 10906 4880 10908
rect 4936 10906 4960 10908
rect 5016 10906 5040 10908
rect 5096 10906 5120 10908
rect 5176 10906 5182 10908
rect 4936 10854 4938 10906
rect 5118 10854 5120 10906
rect 4874 10852 4880 10854
rect 4936 10852 4960 10854
rect 5016 10852 5040 10854
rect 5096 10852 5120 10854
rect 5176 10852 5182 10854
rect 4874 10843 5182 10852
rect 4712 10056 4764 10062
rect 4712 9998 4764 10004
rect 4804 9920 4856 9926
rect 4804 9862 4856 9868
rect 4816 9042 4844 9862
rect 4874 9820 5182 9829
rect 4874 9818 4880 9820
rect 4936 9818 4960 9820
rect 5016 9818 5040 9820
rect 5096 9818 5120 9820
rect 5176 9818 5182 9820
rect 4936 9766 4938 9818
rect 5118 9766 5120 9818
rect 4874 9764 4880 9766
rect 4936 9764 4960 9766
rect 5016 9764 5040 9766
rect 5096 9764 5120 9766
rect 5176 9764 5182 9766
rect 4874 9755 5182 9764
rect 4804 9036 4856 9042
rect 4804 8978 4856 8984
rect 4816 8498 4844 8978
rect 4874 8732 5182 8741
rect 4874 8730 4880 8732
rect 4936 8730 4960 8732
rect 5016 8730 5040 8732
rect 5096 8730 5120 8732
rect 5176 8730 5182 8732
rect 4936 8678 4938 8730
rect 5118 8678 5120 8730
rect 4874 8676 4880 8678
rect 4936 8676 4960 8678
rect 5016 8676 5040 8678
rect 5096 8676 5120 8678
rect 5176 8676 5182 8678
rect 4874 8667 5182 8676
rect 4804 8492 4856 8498
rect 4804 8434 4856 8440
rect 4620 7948 4672 7954
rect 4620 7890 4672 7896
rect 4804 7880 4856 7886
rect 4804 7822 4856 7828
rect 4816 7546 4844 7822
rect 4874 7644 5182 7653
rect 4874 7642 4880 7644
rect 4936 7642 4960 7644
rect 5016 7642 5040 7644
rect 5096 7642 5120 7644
rect 5176 7642 5182 7644
rect 4936 7590 4938 7642
rect 5118 7590 5120 7642
rect 4874 7588 4880 7590
rect 4936 7588 4960 7590
rect 5016 7588 5040 7590
rect 5096 7588 5120 7590
rect 5176 7588 5182 7590
rect 4874 7579 5182 7588
rect 5276 7546 5304 12406
rect 5356 11756 5408 11762
rect 5356 11698 5408 11704
rect 5368 11218 5396 11698
rect 5356 11212 5408 11218
rect 5356 11154 5408 11160
rect 5368 10470 5396 11154
rect 5356 10464 5408 10470
rect 5356 10406 5408 10412
rect 5368 10130 5396 10406
rect 5460 10130 5488 14232
rect 5920 13870 5948 14418
rect 6196 14414 6224 14758
rect 6184 14408 6236 14414
rect 6184 14350 6236 14356
rect 6736 14408 6788 14414
rect 6736 14350 6788 14356
rect 6748 13938 6776 14350
rect 6736 13932 6788 13938
rect 6736 13874 6788 13880
rect 7012 13932 7064 13938
rect 7012 13874 7064 13880
rect 7564 13932 7616 13938
rect 7564 13874 7616 13880
rect 5908 13864 5960 13870
rect 5908 13806 5960 13812
rect 6184 12776 6236 12782
rect 6184 12718 6236 12724
rect 6196 12306 6224 12718
rect 6184 12300 6236 12306
rect 6184 12242 6236 12248
rect 5540 11688 5592 11694
rect 5540 11630 5592 11636
rect 5552 11150 5580 11630
rect 5540 11144 5592 11150
rect 5592 11104 5672 11132
rect 5540 11086 5592 11092
rect 5356 10124 5408 10130
rect 5356 10066 5408 10072
rect 5448 10124 5500 10130
rect 5448 10066 5500 10072
rect 5540 10056 5592 10062
rect 5540 9998 5592 10004
rect 5356 8968 5408 8974
rect 5356 8910 5408 8916
rect 5368 8498 5396 8910
rect 5552 8498 5580 9998
rect 5644 9042 5672 11104
rect 5816 11076 5868 11082
rect 5816 11018 5868 11024
rect 5828 10810 5856 11018
rect 6748 11014 6776 13874
rect 6920 13796 6972 13802
rect 6920 13738 6972 13744
rect 6932 13326 6960 13738
rect 7024 13326 7052 13874
rect 6920 13320 6972 13326
rect 6920 13262 6972 13268
rect 7012 13320 7064 13326
rect 7012 13262 7064 13268
rect 7024 12102 7052 13262
rect 7576 13258 7604 13874
rect 7104 13252 7156 13258
rect 7104 13194 7156 13200
rect 7564 13252 7616 13258
rect 7564 13194 7616 13200
rect 7116 12986 7144 13194
rect 7104 12980 7156 12986
rect 7104 12922 7156 12928
rect 7196 12844 7248 12850
rect 7196 12786 7248 12792
rect 7472 12844 7524 12850
rect 7472 12786 7524 12792
rect 7012 12096 7064 12102
rect 7012 12038 7064 12044
rect 7208 11286 7236 12786
rect 7484 12306 7512 12786
rect 7472 12300 7524 12306
rect 7472 12242 7524 12248
rect 7668 11830 7696 14962
rect 8220 13462 8248 16050
rect 8312 15910 8340 16458
rect 8300 15904 8352 15910
rect 8300 15846 8352 15852
rect 8312 15570 8340 15846
rect 8300 15564 8352 15570
rect 8300 15506 8352 15512
rect 8312 15026 8340 15506
rect 8404 15502 8432 16544
rect 8484 16526 8536 16532
rect 8484 16448 8536 16454
rect 8588 16436 8616 17138
rect 8536 16408 8616 16436
rect 8484 16390 8536 16396
rect 8496 15638 8524 16390
rect 8680 15994 8708 18090
rect 9232 17746 9260 21966
rect 9416 18970 9444 21966
rect 10600 20936 10652 20942
rect 10600 20878 10652 20884
rect 11794 20904 11850 20913
rect 10612 19922 10640 20878
rect 11152 20868 11204 20874
rect 11794 20839 11850 20848
rect 11152 20810 11204 20816
rect 11164 20602 11192 20810
rect 11152 20596 11204 20602
rect 11152 20538 11204 20544
rect 11808 20398 11836 20839
rect 11796 20392 11848 20398
rect 11796 20334 11848 20340
rect 11980 20324 12032 20330
rect 11980 20266 12032 20272
rect 11992 19922 12020 20266
rect 10600 19916 10652 19922
rect 10600 19858 10652 19864
rect 11980 19916 12032 19922
rect 11980 19858 12032 19864
rect 10048 19712 10100 19718
rect 10048 19654 10100 19660
rect 9680 19168 9732 19174
rect 9680 19110 9732 19116
rect 9404 18964 9456 18970
rect 9404 18906 9456 18912
rect 9692 18766 9720 19110
rect 10060 18766 10088 19654
rect 9404 18760 9456 18766
rect 9404 18702 9456 18708
rect 9680 18760 9732 18766
rect 9680 18702 9732 18708
rect 10048 18760 10100 18766
rect 10048 18702 10100 18708
rect 9416 18358 9444 18702
rect 9956 18624 10008 18630
rect 9956 18566 10008 18572
rect 9404 18352 9456 18358
rect 9404 18294 9456 18300
rect 9588 18284 9640 18290
rect 9588 18226 9640 18232
rect 9404 18216 9456 18222
rect 9404 18158 9456 18164
rect 9220 17740 9272 17746
rect 9220 17682 9272 17688
rect 9128 17672 9180 17678
rect 9128 17614 9180 17620
rect 9036 16584 9088 16590
rect 9036 16526 9088 16532
rect 8944 16516 8996 16522
rect 8944 16458 8996 16464
rect 8760 16448 8812 16454
rect 8760 16390 8812 16396
rect 8772 16182 8800 16390
rect 8760 16176 8812 16182
rect 8760 16118 8812 16124
rect 8956 16114 8984 16458
rect 9048 16114 9076 16526
rect 8944 16108 8996 16114
rect 8944 16050 8996 16056
rect 9036 16108 9088 16114
rect 9036 16050 9088 16056
rect 8852 16040 8904 16046
rect 8680 15966 8800 15994
rect 8852 15982 8904 15988
rect 8484 15632 8536 15638
rect 8484 15574 8536 15580
rect 8772 15502 8800 15966
rect 8864 15638 8892 15982
rect 8852 15632 8904 15638
rect 8852 15574 8904 15580
rect 9048 15570 9076 16050
rect 9036 15564 9088 15570
rect 9036 15506 9088 15512
rect 8392 15496 8444 15502
rect 8392 15438 8444 15444
rect 8576 15496 8628 15502
rect 8576 15438 8628 15444
rect 8760 15496 8812 15502
rect 8760 15438 8812 15444
rect 8404 15026 8432 15438
rect 8300 15020 8352 15026
rect 8300 14962 8352 14968
rect 8392 15020 8444 15026
rect 8392 14962 8444 14968
rect 8404 14550 8432 14962
rect 8392 14544 8444 14550
rect 8392 14486 8444 14492
rect 8300 13932 8352 13938
rect 8300 13874 8352 13880
rect 8208 13456 8260 13462
rect 8208 13398 8260 13404
rect 8208 13320 8260 13326
rect 8312 13308 8340 13874
rect 8588 13802 8616 15438
rect 8668 13864 8720 13870
rect 8668 13806 8720 13812
rect 8576 13796 8628 13802
rect 8576 13738 8628 13744
rect 8680 13394 8708 13806
rect 8772 13530 8800 15438
rect 9140 15434 9168 17614
rect 9416 17542 9444 18158
rect 9496 18148 9548 18154
rect 9496 18090 9548 18096
rect 9508 17678 9536 18090
rect 9600 17746 9628 18226
rect 9864 18080 9916 18086
rect 9864 18022 9916 18028
rect 9876 17814 9904 18022
rect 9864 17808 9916 17814
rect 9864 17750 9916 17756
rect 9588 17740 9640 17746
rect 9588 17682 9640 17688
rect 9496 17672 9548 17678
rect 9496 17614 9548 17620
rect 9404 17536 9456 17542
rect 9404 17478 9456 17484
rect 9416 16794 9444 17478
rect 9876 17202 9904 17750
rect 9968 17202 9996 18566
rect 10060 18290 10088 18702
rect 10324 18624 10376 18630
rect 10324 18566 10376 18572
rect 10048 18284 10100 18290
rect 10048 18226 10100 18232
rect 10336 17678 10364 18566
rect 10324 17672 10376 17678
rect 10324 17614 10376 17620
rect 10612 17270 10640 19858
rect 10968 18896 11020 18902
rect 10968 18838 11020 18844
rect 10980 17678 11008 18838
rect 11060 18284 11112 18290
rect 11060 18226 11112 18232
rect 11072 17882 11100 18226
rect 11888 18148 11940 18154
rect 11888 18090 11940 18096
rect 11060 17876 11112 17882
rect 11060 17818 11112 17824
rect 10968 17672 11020 17678
rect 10968 17614 11020 17620
rect 10784 17536 10836 17542
rect 10784 17478 10836 17484
rect 11796 17536 11848 17542
rect 11796 17478 11848 17484
rect 10600 17264 10652 17270
rect 10600 17206 10652 17212
rect 10796 17202 10824 17478
rect 11808 17202 11836 17478
rect 11900 17202 11928 18090
rect 11992 17678 12020 19858
rect 12072 18216 12124 18222
rect 12072 18158 12124 18164
rect 11980 17672 12032 17678
rect 11980 17614 12032 17620
rect 9864 17196 9916 17202
rect 9864 17138 9916 17144
rect 9956 17196 10008 17202
rect 9956 17138 10008 17144
rect 10784 17196 10836 17202
rect 10784 17138 10836 17144
rect 11796 17196 11848 17202
rect 11796 17138 11848 17144
rect 11888 17196 11940 17202
rect 11888 17138 11940 17144
rect 11980 17196 12032 17202
rect 12084 17184 12112 18158
rect 12176 17746 12204 23462
rect 12268 23118 12296 23666
rect 12544 23118 12572 23820
rect 12256 23112 12308 23118
rect 12256 23054 12308 23060
rect 12532 23112 12584 23118
rect 12532 23054 12584 23060
rect 12624 23112 12676 23118
rect 12624 23054 12676 23060
rect 12636 22438 12664 23054
rect 12728 22506 12756 24142
rect 12912 23118 12940 25094
rect 13004 24206 13032 26182
rect 13096 25362 13124 26318
rect 13176 26240 13228 26246
rect 13176 26182 13228 26188
rect 13188 25906 13216 26182
rect 13176 25900 13228 25906
rect 13176 25842 13228 25848
rect 20088 25702 20116 27610
rect 20260 27464 20312 27470
rect 20260 27406 20312 27412
rect 20168 27396 20220 27402
rect 20168 27338 20220 27344
rect 20180 26790 20208 27338
rect 20272 26994 20300 27406
rect 20364 27130 20392 28018
rect 21088 28008 21140 28014
rect 21088 27950 21140 27956
rect 20996 27940 21048 27946
rect 20996 27882 21048 27888
rect 20812 27668 20864 27674
rect 20812 27610 20864 27616
rect 20824 27334 20852 27610
rect 20904 27464 20956 27470
rect 20904 27406 20956 27412
rect 20812 27328 20864 27334
rect 20812 27270 20864 27276
rect 20352 27124 20404 27130
rect 20352 27066 20404 27072
rect 20626 27024 20682 27033
rect 20260 26988 20312 26994
rect 20312 26948 20392 26976
rect 20626 26959 20628 26968
rect 20260 26930 20312 26936
rect 20168 26784 20220 26790
rect 20168 26726 20220 26732
rect 20180 26586 20208 26726
rect 20168 26580 20220 26586
rect 20168 26522 20220 26528
rect 20180 26382 20208 26522
rect 20364 26382 20392 26948
rect 20680 26959 20682 26968
rect 20628 26930 20680 26936
rect 20444 26920 20496 26926
rect 20444 26862 20496 26868
rect 20456 26790 20484 26862
rect 20628 26852 20680 26858
rect 20628 26794 20680 26800
rect 20444 26784 20496 26790
rect 20444 26726 20496 26732
rect 20640 26450 20668 26794
rect 20628 26444 20680 26450
rect 20628 26386 20680 26392
rect 20824 26382 20852 27270
rect 20916 27062 20944 27406
rect 21008 27402 21036 27882
rect 21100 27606 21128 27950
rect 21376 27674 21404 28494
rect 21456 28484 21508 28490
rect 21456 28426 21508 28432
rect 21364 27668 21416 27674
rect 21364 27610 21416 27616
rect 21468 27606 21496 28426
rect 21640 28076 21692 28082
rect 22100 28076 22152 28082
rect 21640 28018 21692 28024
rect 21928 28036 22100 28064
rect 21548 27872 21600 27878
rect 21548 27814 21600 27820
rect 21088 27600 21140 27606
rect 21088 27542 21140 27548
rect 21456 27600 21508 27606
rect 21456 27542 21508 27548
rect 20996 27396 21048 27402
rect 20996 27338 21048 27344
rect 21008 27130 21036 27338
rect 21560 27130 21588 27814
rect 21652 27538 21680 28018
rect 21640 27532 21692 27538
rect 21640 27474 21692 27480
rect 20996 27124 21048 27130
rect 20996 27066 21048 27072
rect 21548 27124 21600 27130
rect 21548 27066 21600 27072
rect 21928 27062 21956 28036
rect 22100 28018 22152 28024
rect 22100 27872 22152 27878
rect 22100 27814 22152 27820
rect 22112 27538 22140 27814
rect 22296 27674 22324 28494
rect 22376 28008 22428 28014
rect 22376 27950 22428 27956
rect 22284 27668 22336 27674
rect 22284 27610 22336 27616
rect 22100 27532 22152 27538
rect 22100 27474 22152 27480
rect 22388 27418 22416 27950
rect 22560 27600 22612 27606
rect 22560 27542 22612 27548
rect 22192 27396 22244 27402
rect 22388 27390 22508 27418
rect 22572 27402 22600 27542
rect 22192 27338 22244 27344
rect 20904 27056 20956 27062
rect 20904 26998 20956 27004
rect 21916 27056 21968 27062
rect 21916 26998 21968 27004
rect 20996 26988 21048 26994
rect 20996 26930 21048 26936
rect 21456 26988 21508 26994
rect 21456 26930 21508 26936
rect 20168 26376 20220 26382
rect 20168 26318 20220 26324
rect 20352 26376 20404 26382
rect 20352 26318 20404 26324
rect 20812 26376 20864 26382
rect 20812 26318 20864 26324
rect 20628 26308 20680 26314
rect 20628 26250 20680 26256
rect 20076 25696 20128 25702
rect 20076 25638 20128 25644
rect 20444 25696 20496 25702
rect 20444 25638 20496 25644
rect 20456 25498 20484 25638
rect 20640 25498 20668 26250
rect 20824 26246 20852 26318
rect 20812 26240 20864 26246
rect 20812 26182 20864 26188
rect 20444 25492 20496 25498
rect 20444 25434 20496 25440
rect 20628 25492 20680 25498
rect 20628 25434 20680 25440
rect 15568 25424 15620 25430
rect 15568 25366 15620 25372
rect 13084 25356 13136 25362
rect 13084 25298 13136 25304
rect 15292 25356 15344 25362
rect 15292 25298 15344 25304
rect 13096 24886 13124 25298
rect 15200 25220 15252 25226
rect 15200 25162 15252 25168
rect 13084 24880 13136 24886
rect 13084 24822 13136 24828
rect 13360 24880 13412 24886
rect 13360 24822 13412 24828
rect 13176 24812 13228 24818
rect 13176 24754 13228 24760
rect 13084 24608 13136 24614
rect 13084 24550 13136 24556
rect 12992 24200 13044 24206
rect 12992 24142 13044 24148
rect 12992 23520 13044 23526
rect 12992 23462 13044 23468
rect 13004 23322 13032 23462
rect 12992 23316 13044 23322
rect 12992 23258 13044 23264
rect 12900 23112 12952 23118
rect 12900 23054 12952 23060
rect 13096 22574 13124 24550
rect 13188 24410 13216 24754
rect 13176 24404 13228 24410
rect 13176 24346 13228 24352
rect 13372 24206 13400 24822
rect 15212 24818 15240 25162
rect 15304 24818 15332 25298
rect 15580 25294 15608 25366
rect 15568 25288 15620 25294
rect 15568 25230 15620 25236
rect 16120 25288 16172 25294
rect 16120 25230 16172 25236
rect 15580 24818 15608 25230
rect 14096 24812 14148 24818
rect 14096 24754 14148 24760
rect 15200 24812 15252 24818
rect 15200 24754 15252 24760
rect 15292 24812 15344 24818
rect 15292 24754 15344 24760
rect 15568 24812 15620 24818
rect 15568 24754 15620 24760
rect 14108 24206 14136 24754
rect 15580 24682 15608 24754
rect 16132 24750 16160 25230
rect 20824 25226 20852 26182
rect 21008 25498 21036 26930
rect 21468 26518 21496 26930
rect 22204 26874 22232 27338
rect 22480 27062 22508 27390
rect 22560 27396 22612 27402
rect 22560 27338 22612 27344
rect 22664 27130 22692 28494
rect 23020 27464 23072 27470
rect 23020 27406 23072 27412
rect 23112 27464 23164 27470
rect 23112 27406 23164 27412
rect 22928 27328 22980 27334
rect 22928 27270 22980 27276
rect 22652 27124 22704 27130
rect 22652 27066 22704 27072
rect 22284 27056 22336 27062
rect 22282 27024 22284 27033
rect 22468 27056 22520 27062
rect 22336 27024 22338 27033
rect 22338 26982 22416 27010
rect 22468 26998 22520 27004
rect 22282 26959 22338 26968
rect 22204 26858 22324 26874
rect 21824 26852 21876 26858
rect 22204 26852 22336 26858
rect 22204 26846 22284 26852
rect 21824 26794 21876 26800
rect 22284 26794 22336 26800
rect 21456 26512 21508 26518
rect 21456 26454 21508 26460
rect 21836 26382 21864 26794
rect 21824 26376 21876 26382
rect 21824 26318 21876 26324
rect 21836 25906 21864 26318
rect 21824 25900 21876 25906
rect 21824 25842 21876 25848
rect 20996 25492 21048 25498
rect 20996 25434 21048 25440
rect 16672 25220 16724 25226
rect 16672 25162 16724 25168
rect 20812 25220 20864 25226
rect 20812 25162 20864 25168
rect 16684 24954 16712 25162
rect 21008 25158 21036 25434
rect 22388 25362 22416 26982
rect 22480 26314 22508 26998
rect 22940 26994 22968 27270
rect 23032 26994 23060 27406
rect 23124 27062 23152 27406
rect 23308 27130 23336 28494
rect 23388 28076 23440 28082
rect 23388 28018 23440 28024
rect 23400 27470 23428 28018
rect 23952 27674 23980 28494
rect 24032 27940 24084 27946
rect 24032 27882 24084 27888
rect 23940 27668 23992 27674
rect 23940 27610 23992 27616
rect 24044 27470 24072 27882
rect 24596 27674 24624 28494
rect 24964 28218 24992 28494
rect 24952 28212 25004 28218
rect 24952 28154 25004 28160
rect 24952 28076 25004 28082
rect 24952 28018 25004 28024
rect 25044 28076 25096 28082
rect 25044 28018 25096 28024
rect 24584 27668 24636 27674
rect 24584 27610 24636 27616
rect 24676 27668 24728 27674
rect 24676 27610 24728 27616
rect 24688 27554 24716 27610
rect 24596 27526 24716 27554
rect 24860 27532 24912 27538
rect 23388 27464 23440 27470
rect 23388 27406 23440 27412
rect 24032 27464 24084 27470
rect 24032 27406 24084 27412
rect 24216 27464 24268 27470
rect 24216 27406 24268 27412
rect 24400 27464 24452 27470
rect 24400 27406 24452 27412
rect 23756 27396 23808 27402
rect 23756 27338 23808 27344
rect 23296 27124 23348 27130
rect 23296 27066 23348 27072
rect 23112 27056 23164 27062
rect 23112 26998 23164 27004
rect 22652 26988 22704 26994
rect 22652 26930 22704 26936
rect 22928 26988 22980 26994
rect 22928 26930 22980 26936
rect 23020 26988 23072 26994
rect 23020 26930 23072 26936
rect 23664 26988 23716 26994
rect 23664 26930 23716 26936
rect 22664 26586 22692 26930
rect 22652 26580 22704 26586
rect 22652 26522 22704 26528
rect 23676 26314 23704 26930
rect 22468 26308 22520 26314
rect 22468 26250 22520 26256
rect 23020 26308 23072 26314
rect 23020 26250 23072 26256
rect 23664 26308 23716 26314
rect 23664 26250 23716 26256
rect 22376 25356 22428 25362
rect 22376 25298 22428 25304
rect 21824 25288 21876 25294
rect 21824 25230 21876 25236
rect 16764 25152 16816 25158
rect 16764 25094 16816 25100
rect 20996 25152 21048 25158
rect 20996 25094 21048 25100
rect 16672 24948 16724 24954
rect 16672 24890 16724 24896
rect 16684 24818 16712 24890
rect 16776 24818 16804 25094
rect 16304 24812 16356 24818
rect 16304 24754 16356 24760
rect 16580 24812 16632 24818
rect 16580 24754 16632 24760
rect 16672 24812 16724 24818
rect 16672 24754 16724 24760
rect 16764 24812 16816 24818
rect 16764 24754 16816 24760
rect 20628 24812 20680 24818
rect 20628 24754 20680 24760
rect 21732 24812 21784 24818
rect 21732 24754 21784 24760
rect 16120 24744 16172 24750
rect 16120 24686 16172 24692
rect 15568 24676 15620 24682
rect 15568 24618 15620 24624
rect 15752 24608 15804 24614
rect 15752 24550 15804 24556
rect 15936 24608 15988 24614
rect 15936 24550 15988 24556
rect 13360 24200 13412 24206
rect 13360 24142 13412 24148
rect 14096 24200 14148 24206
rect 14096 24142 14148 24148
rect 13372 23798 13400 24142
rect 14556 24132 14608 24138
rect 14556 24074 14608 24080
rect 15568 24132 15620 24138
rect 15568 24074 15620 24080
rect 13360 23792 13412 23798
rect 13360 23734 13412 23740
rect 14568 23730 14596 24074
rect 14556 23724 14608 23730
rect 14556 23666 14608 23672
rect 14280 23180 14332 23186
rect 14280 23122 14332 23128
rect 13268 23112 13320 23118
rect 13268 23054 13320 23060
rect 13544 23112 13596 23118
rect 13544 23054 13596 23060
rect 13084 22568 13136 22574
rect 13084 22510 13136 22516
rect 13280 22506 13308 23054
rect 13556 22778 13584 23054
rect 14096 22976 14148 22982
rect 14096 22918 14148 22924
rect 13544 22772 13596 22778
rect 13544 22714 13596 22720
rect 14108 22710 14136 22918
rect 14096 22704 14148 22710
rect 14096 22646 14148 22652
rect 13360 22636 13412 22642
rect 13360 22578 13412 22584
rect 12716 22500 12768 22506
rect 12716 22442 12768 22448
rect 13268 22500 13320 22506
rect 13268 22442 13320 22448
rect 12624 22432 12676 22438
rect 12624 22374 12676 22380
rect 12808 22432 12860 22438
rect 12808 22374 12860 22380
rect 12348 22024 12400 22030
rect 12348 21966 12400 21972
rect 12360 21554 12388 21966
rect 12348 21548 12400 21554
rect 12348 21490 12400 21496
rect 12360 21146 12388 21490
rect 12532 21412 12584 21418
rect 12532 21354 12584 21360
rect 12348 21140 12400 21146
rect 12348 21082 12400 21088
rect 12256 20868 12308 20874
rect 12256 20810 12308 20816
rect 12268 19786 12296 20810
rect 12544 20806 12572 21354
rect 12716 21140 12768 21146
rect 12716 21082 12768 21088
rect 12532 20800 12584 20806
rect 12530 20768 12532 20777
rect 12624 20800 12676 20806
rect 12584 20768 12586 20777
rect 12624 20742 12676 20748
rect 12530 20703 12586 20712
rect 12532 20528 12584 20534
rect 12530 20496 12532 20505
rect 12584 20496 12586 20505
rect 12530 20431 12586 20440
rect 12348 20392 12400 20398
rect 12348 20334 12400 20340
rect 12360 20058 12388 20334
rect 12440 20324 12492 20330
rect 12440 20266 12492 20272
rect 12348 20052 12400 20058
rect 12348 19994 12400 20000
rect 12256 19780 12308 19786
rect 12256 19722 12308 19728
rect 12268 19514 12296 19722
rect 12256 19508 12308 19514
rect 12256 19450 12308 19456
rect 12452 18290 12480 20266
rect 12636 19922 12664 20742
rect 12728 20602 12756 21082
rect 12716 20596 12768 20602
rect 12716 20538 12768 20544
rect 12716 20460 12768 20466
rect 12716 20402 12768 20408
rect 12728 19922 12756 20402
rect 12820 20398 12848 22374
rect 13084 21684 13136 21690
rect 13084 21626 13136 21632
rect 12898 21584 12954 21593
rect 13096 21554 13124 21626
rect 12898 21519 12900 21528
rect 12952 21519 12954 21528
rect 13084 21548 13136 21554
rect 12900 21490 12952 21496
rect 13084 21490 13136 21496
rect 13176 21548 13228 21554
rect 13176 21490 13228 21496
rect 13096 21418 13124 21490
rect 13188 21418 13216 21490
rect 13084 21412 13136 21418
rect 13084 21354 13136 21360
rect 13176 21412 13228 21418
rect 13176 21354 13228 21360
rect 12992 21344 13044 21350
rect 12992 21286 13044 21292
rect 13004 21010 13032 21286
rect 12992 21004 13044 21010
rect 12992 20946 13044 20952
rect 13084 20936 13136 20942
rect 13084 20878 13136 20884
rect 12992 20868 13044 20874
rect 12992 20810 13044 20816
rect 12808 20392 12860 20398
rect 12808 20334 12860 20340
rect 12808 20256 12860 20262
rect 12808 20198 12860 20204
rect 12624 19916 12676 19922
rect 12624 19858 12676 19864
rect 12716 19916 12768 19922
rect 12716 19858 12768 19864
rect 12440 18284 12492 18290
rect 12440 18226 12492 18232
rect 12636 18222 12664 19858
rect 12728 18426 12756 19858
rect 12716 18420 12768 18426
rect 12716 18362 12768 18368
rect 12624 18216 12676 18222
rect 12624 18158 12676 18164
rect 12624 18080 12676 18086
rect 12624 18022 12676 18028
rect 12164 17740 12216 17746
rect 12164 17682 12216 17688
rect 12032 17156 12112 17184
rect 11980 17138 12032 17144
rect 10876 17128 10928 17134
rect 10876 17070 10928 17076
rect 9772 16992 9824 16998
rect 9772 16934 9824 16940
rect 9404 16788 9456 16794
rect 9404 16730 9456 16736
rect 9784 16658 9812 16934
rect 10888 16726 10916 17070
rect 10876 16720 10928 16726
rect 10876 16662 10928 16668
rect 9772 16652 9824 16658
rect 9772 16594 9824 16600
rect 9784 16114 9812 16594
rect 11152 16448 11204 16454
rect 11152 16390 11204 16396
rect 9772 16108 9824 16114
rect 9772 16050 9824 16056
rect 9864 15496 9916 15502
rect 9864 15438 9916 15444
rect 9128 15428 9180 15434
rect 9128 15370 9180 15376
rect 9876 15094 9904 15438
rect 9864 15088 9916 15094
rect 9864 15030 9916 15036
rect 10232 15088 10284 15094
rect 10232 15030 10284 15036
rect 9588 13932 9640 13938
rect 9588 13874 9640 13880
rect 9680 13932 9732 13938
rect 9680 13874 9732 13880
rect 9128 13728 9180 13734
rect 9128 13670 9180 13676
rect 9220 13728 9272 13734
rect 9220 13670 9272 13676
rect 8760 13524 8812 13530
rect 8760 13466 8812 13472
rect 9140 13394 9168 13670
rect 8668 13388 8720 13394
rect 8668 13330 8720 13336
rect 9128 13388 9180 13394
rect 9128 13330 9180 13336
rect 9232 13326 9260 13670
rect 8260 13280 8340 13308
rect 8208 13262 8260 13268
rect 8312 12986 8340 13280
rect 8484 13320 8536 13326
rect 8484 13262 8536 13268
rect 9220 13320 9272 13326
rect 9220 13262 9272 13268
rect 8300 12980 8352 12986
rect 8300 12922 8352 12928
rect 8496 12850 8524 13262
rect 9600 12850 9628 13874
rect 9692 13258 9720 13874
rect 10244 13530 10272 15030
rect 11164 14414 11192 16390
rect 11520 15020 11572 15026
rect 11520 14962 11572 14968
rect 11704 15020 11756 15026
rect 11704 14962 11756 14968
rect 11888 15020 11940 15026
rect 11888 14962 11940 14968
rect 11152 14408 11204 14414
rect 11152 14350 11204 14356
rect 11244 14408 11296 14414
rect 11244 14350 11296 14356
rect 10232 13524 10284 13530
rect 10232 13466 10284 13472
rect 10416 13524 10468 13530
rect 10416 13466 10468 13472
rect 10232 13320 10284 13326
rect 10232 13262 10284 13268
rect 9680 13252 9732 13258
rect 9680 13194 9732 13200
rect 8484 12844 8536 12850
rect 8484 12786 8536 12792
rect 9588 12844 9640 12850
rect 9588 12786 9640 12792
rect 9692 12782 9720 13194
rect 10048 13184 10100 13190
rect 10048 13126 10100 13132
rect 10060 13025 10088 13126
rect 10046 13016 10102 13025
rect 10046 12951 10102 12960
rect 9680 12776 9732 12782
rect 9680 12718 9732 12724
rect 8484 12232 8536 12238
rect 8484 12174 8536 12180
rect 7656 11824 7708 11830
rect 7656 11766 7708 11772
rect 7196 11280 7248 11286
rect 7196 11222 7248 11228
rect 7564 11212 7616 11218
rect 7564 11154 7616 11160
rect 6460 11008 6512 11014
rect 6460 10950 6512 10956
rect 6736 11008 6788 11014
rect 6736 10950 6788 10956
rect 5816 10804 5868 10810
rect 5816 10746 5868 10752
rect 6472 10742 6500 10950
rect 6460 10736 6512 10742
rect 6460 10678 6512 10684
rect 6368 10668 6420 10674
rect 6288 10628 6368 10656
rect 6288 9178 6316 10628
rect 6368 10610 6420 10616
rect 6472 10606 6500 10678
rect 6460 10600 6512 10606
rect 6460 10542 6512 10548
rect 6748 10062 6776 10950
rect 7576 10606 7604 11154
rect 8496 10742 8524 12174
rect 8760 11756 8812 11762
rect 8760 11698 8812 11704
rect 8772 11626 8800 11698
rect 9220 11688 9272 11694
rect 9220 11630 9272 11636
rect 8760 11620 8812 11626
rect 8760 11562 8812 11568
rect 8576 11144 8628 11150
rect 8772 11098 8800 11562
rect 8628 11092 8800 11098
rect 8576 11086 8800 11092
rect 8588 11070 8800 11086
rect 8484 10736 8536 10742
rect 8484 10678 8536 10684
rect 7564 10600 7616 10606
rect 7564 10542 7616 10548
rect 8392 10600 8444 10606
rect 8392 10542 8444 10548
rect 8404 10266 8432 10542
rect 8392 10260 8444 10266
rect 8392 10202 8444 10208
rect 8300 10192 8352 10198
rect 8352 10140 8432 10146
rect 8300 10134 8432 10140
rect 8312 10118 8432 10134
rect 8404 10062 8432 10118
rect 6736 10056 6788 10062
rect 6736 9998 6788 10004
rect 8392 10056 8444 10062
rect 8392 9998 8444 10004
rect 8300 9988 8352 9994
rect 8300 9930 8352 9936
rect 6276 9172 6328 9178
rect 6276 9114 6328 9120
rect 5632 9036 5684 9042
rect 5632 8978 5684 8984
rect 5816 8968 5868 8974
rect 5816 8910 5868 8916
rect 5908 8968 5960 8974
rect 6092 8968 6144 8974
rect 5908 8910 5960 8916
rect 6012 8928 6092 8956
rect 5828 8634 5856 8910
rect 5920 8838 5948 8910
rect 5908 8832 5960 8838
rect 5908 8774 5960 8780
rect 5816 8628 5868 8634
rect 5816 8570 5868 8576
rect 5356 8492 5408 8498
rect 5356 8434 5408 8440
rect 5540 8492 5592 8498
rect 5540 8434 5592 8440
rect 5816 8492 5868 8498
rect 5816 8434 5868 8440
rect 5368 8090 5396 8434
rect 5356 8084 5408 8090
rect 5356 8026 5408 8032
rect 5448 7880 5500 7886
rect 5448 7822 5500 7828
rect 4804 7540 4856 7546
rect 4804 7482 4856 7488
rect 5264 7540 5316 7546
rect 5264 7482 5316 7488
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 5276 6934 5304 7482
rect 5460 7342 5488 7822
rect 5552 7410 5580 8434
rect 5828 8294 5856 8434
rect 5920 8430 5948 8774
rect 6012 8498 6040 8928
rect 6092 8910 6144 8916
rect 8116 8968 8168 8974
rect 8116 8910 8168 8916
rect 6184 8900 6236 8906
rect 6184 8842 6236 8848
rect 8024 8900 8076 8906
rect 8024 8842 8076 8848
rect 6196 8498 6224 8842
rect 8036 8498 8064 8842
rect 6000 8492 6052 8498
rect 6000 8434 6052 8440
rect 6184 8492 6236 8498
rect 6184 8434 6236 8440
rect 8024 8492 8076 8498
rect 8024 8434 8076 8440
rect 5908 8424 5960 8430
rect 5908 8366 5960 8372
rect 5816 8288 5868 8294
rect 5816 8230 5868 8236
rect 5828 7954 5856 8230
rect 6552 8084 6604 8090
rect 6552 8026 6604 8032
rect 5816 7948 5868 7954
rect 5816 7890 5868 7896
rect 5828 7410 5856 7890
rect 6092 7880 6144 7886
rect 6092 7822 6144 7828
rect 5540 7404 5592 7410
rect 5540 7346 5592 7352
rect 5816 7404 5868 7410
rect 5816 7346 5868 7352
rect 5448 7336 5500 7342
rect 5448 7278 5500 7284
rect 5540 7200 5592 7206
rect 5540 7142 5592 7148
rect 5264 6928 5316 6934
rect 5264 6870 5316 6876
rect 5552 6866 5580 7142
rect 5540 6860 5592 6866
rect 5540 6802 5592 6808
rect 6000 6656 6052 6662
rect 6000 6598 6052 6604
rect 4874 6556 5182 6565
rect 4874 6554 4880 6556
rect 4936 6554 4960 6556
rect 5016 6554 5040 6556
rect 5096 6554 5120 6556
rect 5176 6554 5182 6556
rect 4936 6502 4938 6554
rect 5118 6502 5120 6554
rect 4874 6500 4880 6502
rect 4936 6500 4960 6502
rect 5016 6500 5040 6502
rect 5096 6500 5120 6502
rect 5176 6500 5182 6502
rect 4874 6491 5182 6500
rect 6012 6322 6040 6598
rect 6000 6316 6052 6322
rect 6000 6258 6052 6264
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4874 5468 5182 5477
rect 4874 5466 4880 5468
rect 4936 5466 4960 5468
rect 5016 5466 5040 5468
rect 5096 5466 5120 5468
rect 5176 5466 5182 5468
rect 4936 5414 4938 5466
rect 5118 5414 5120 5466
rect 4874 5412 4880 5414
rect 4936 5412 4960 5414
rect 5016 5412 5040 5414
rect 5096 5412 5120 5414
rect 5176 5412 5182 5414
rect 4874 5403 5182 5412
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4874 4380 5182 4389
rect 4874 4378 4880 4380
rect 4936 4378 4960 4380
rect 5016 4378 5040 4380
rect 5096 4378 5120 4380
rect 5176 4378 5182 4380
rect 4936 4326 4938 4378
rect 5118 4326 5120 4378
rect 4874 4324 4880 4326
rect 4936 4324 4960 4326
rect 5016 4324 5040 4326
rect 5096 4324 5120 4326
rect 5176 4324 5182 4326
rect 4874 4315 5182 4324
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4874 3292 5182 3301
rect 4874 3290 4880 3292
rect 4936 3290 4960 3292
rect 5016 3290 5040 3292
rect 5096 3290 5120 3292
rect 5176 3290 5182 3292
rect 4936 3238 4938 3290
rect 5118 3238 5120 3290
rect 4874 3236 4880 3238
rect 4936 3236 4960 3238
rect 5016 3236 5040 3238
rect 5096 3236 5120 3238
rect 5176 3236 5182 3238
rect 4874 3227 5182 3236
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 6104 2650 6132 7822
rect 6564 7410 6592 8026
rect 8036 7546 8064 8434
rect 8128 8430 8156 8910
rect 8116 8424 8168 8430
rect 8116 8366 8168 8372
rect 8312 7546 8340 9930
rect 8496 8090 8524 10678
rect 8588 10674 8616 11070
rect 8668 11008 8720 11014
rect 8668 10950 8720 10956
rect 8680 10810 8708 10950
rect 8668 10804 8720 10810
rect 8668 10746 8720 10752
rect 8576 10668 8628 10674
rect 8576 10610 8628 10616
rect 8484 8084 8536 8090
rect 8484 8026 8536 8032
rect 8024 7540 8076 7546
rect 8024 7482 8076 7488
rect 8300 7540 8352 7546
rect 8300 7482 8352 7488
rect 8496 7410 8524 8026
rect 8588 7410 8616 10610
rect 8680 10266 8708 10746
rect 9232 10674 9260 11630
rect 9588 11552 9640 11558
rect 9588 11494 9640 11500
rect 9600 11150 9628 11494
rect 9588 11144 9640 11150
rect 9588 11086 9640 11092
rect 9220 10668 9272 10674
rect 9220 10610 9272 10616
rect 8852 10532 8904 10538
rect 8852 10474 8904 10480
rect 8668 10260 8720 10266
rect 8668 10202 8720 10208
rect 8864 10130 8892 10474
rect 8852 10124 8904 10130
rect 8852 10066 8904 10072
rect 8760 9920 8812 9926
rect 8760 9862 8812 9868
rect 6552 7404 6604 7410
rect 6552 7346 6604 7352
rect 8024 7404 8076 7410
rect 8024 7346 8076 7352
rect 8392 7404 8444 7410
rect 8392 7346 8444 7352
rect 8484 7404 8536 7410
rect 8484 7346 8536 7352
rect 8576 7404 8628 7410
rect 8576 7346 8628 7352
rect 6564 7206 6592 7346
rect 7564 7268 7616 7274
rect 7564 7210 7616 7216
rect 6552 7200 6604 7206
rect 6552 7142 6604 7148
rect 7576 6934 7604 7210
rect 8036 7002 8064 7346
rect 8024 6996 8076 7002
rect 8024 6938 8076 6944
rect 7564 6928 7616 6934
rect 7564 6870 7616 6876
rect 7576 6798 7604 6870
rect 8404 6866 8432 7346
rect 8496 6934 8524 7346
rect 8484 6928 8536 6934
rect 8484 6870 8536 6876
rect 8392 6860 8444 6866
rect 8392 6802 8444 6808
rect 7564 6792 7616 6798
rect 7564 6734 7616 6740
rect 8404 6662 8432 6802
rect 8772 6798 8800 9862
rect 8864 9654 8892 10066
rect 9692 10062 9720 12718
rect 10244 11762 10272 13262
rect 9864 11756 9916 11762
rect 9864 11698 9916 11704
rect 10232 11756 10284 11762
rect 10232 11698 10284 11704
rect 9772 11688 9824 11694
rect 9772 11630 9824 11636
rect 9784 11150 9812 11630
rect 9772 11144 9824 11150
rect 9772 11086 9824 11092
rect 9876 10810 9904 11698
rect 9956 11144 10008 11150
rect 9956 11086 10008 11092
rect 9864 10804 9916 10810
rect 9864 10746 9916 10752
rect 9772 10736 9824 10742
rect 9772 10678 9824 10684
rect 9036 10056 9088 10062
rect 8956 10016 9036 10044
rect 8852 9648 8904 9654
rect 8852 9590 8904 9596
rect 8956 9382 8984 10016
rect 9036 9998 9088 10004
rect 9496 10056 9548 10062
rect 9496 9998 9548 10004
rect 9680 10056 9732 10062
rect 9680 9998 9732 10004
rect 9508 9654 9536 9998
rect 9588 9988 9640 9994
rect 9588 9930 9640 9936
rect 9600 9722 9628 9930
rect 9588 9716 9640 9722
rect 9588 9658 9640 9664
rect 9496 9648 9548 9654
rect 9496 9590 9548 9596
rect 8944 9376 8996 9382
rect 8944 9318 8996 9324
rect 8956 9178 8984 9318
rect 9508 9194 9536 9590
rect 8944 9172 8996 9178
rect 9508 9166 9628 9194
rect 8944 9114 8996 9120
rect 9600 8906 9628 9166
rect 9680 8968 9732 8974
rect 9680 8910 9732 8916
rect 9588 8900 9640 8906
rect 9588 8842 9640 8848
rect 9600 8566 9628 8842
rect 9692 8634 9720 8910
rect 9680 8628 9732 8634
rect 9680 8570 9732 8576
rect 9588 8560 9640 8566
rect 9588 8502 9640 8508
rect 9588 8424 9640 8430
rect 9588 8366 9640 8372
rect 9600 8090 9628 8366
rect 9588 8084 9640 8090
rect 9588 8026 9640 8032
rect 9128 7880 9180 7886
rect 9128 7822 9180 7828
rect 9588 7880 9640 7886
rect 9588 7822 9640 7828
rect 8852 7540 8904 7546
rect 8852 7482 8904 7488
rect 8864 6798 8892 7482
rect 9140 7410 9168 7822
rect 9036 7404 9088 7410
rect 9036 7346 9088 7352
rect 9128 7404 9180 7410
rect 9128 7346 9180 7352
rect 9048 7206 9076 7346
rect 9036 7200 9088 7206
rect 9036 7142 9088 7148
rect 8576 6792 8628 6798
rect 8576 6734 8628 6740
rect 8760 6792 8812 6798
rect 8760 6734 8812 6740
rect 8852 6792 8904 6798
rect 8852 6734 8904 6740
rect 8484 6724 8536 6730
rect 8484 6666 8536 6672
rect 8392 6656 8444 6662
rect 8392 6598 8444 6604
rect 8392 6248 8444 6254
rect 8392 6190 8444 6196
rect 8404 5710 8432 6190
rect 8496 5914 8524 6666
rect 8588 6322 8616 6734
rect 8668 6656 8720 6662
rect 8668 6598 8720 6604
rect 8576 6316 8628 6322
rect 8576 6258 8628 6264
rect 8484 5908 8536 5914
rect 8484 5850 8536 5856
rect 8680 5710 8708 6598
rect 8772 6186 8800 6734
rect 8944 6316 8996 6322
rect 8944 6258 8996 6264
rect 8760 6180 8812 6186
rect 8760 6122 8812 6128
rect 8956 5778 8984 6258
rect 8944 5772 8996 5778
rect 8944 5714 8996 5720
rect 8392 5704 8444 5710
rect 8392 5646 8444 5652
rect 8668 5704 8720 5710
rect 8668 5646 8720 5652
rect 9048 2774 9076 7142
rect 9140 7002 9168 7346
rect 9600 7342 9628 7822
rect 9784 7546 9812 10678
rect 9864 10668 9916 10674
rect 9968 10656 9996 11086
rect 10428 10674 10456 13466
rect 10968 12776 11020 12782
rect 10968 12718 11020 12724
rect 10980 11830 11008 12718
rect 11164 12442 11192 14350
rect 11256 13938 11284 14350
rect 11244 13932 11296 13938
rect 11244 13874 11296 13880
rect 11152 12436 11204 12442
rect 11152 12378 11204 12384
rect 10968 11824 11020 11830
rect 10968 11766 11020 11772
rect 11060 11824 11112 11830
rect 11060 11766 11112 11772
rect 11072 11354 11100 11766
rect 11334 11656 11390 11665
rect 11334 11591 11336 11600
rect 11388 11591 11390 11600
rect 11336 11562 11388 11568
rect 11152 11552 11204 11558
rect 11152 11494 11204 11500
rect 11060 11348 11112 11354
rect 11060 11290 11112 11296
rect 10600 11144 10652 11150
rect 10600 11086 10652 11092
rect 9916 10628 9996 10656
rect 10416 10668 10468 10674
rect 9864 10610 9916 10616
rect 10416 10610 10468 10616
rect 10428 10470 10456 10610
rect 10416 10464 10468 10470
rect 10416 10406 10468 10412
rect 10612 9042 10640 11086
rect 10692 11076 10744 11082
rect 10692 11018 10744 11024
rect 10876 11076 10928 11082
rect 10876 11018 10928 11024
rect 10704 10538 10732 11018
rect 10692 10532 10744 10538
rect 10692 10474 10744 10480
rect 10600 9036 10652 9042
rect 10600 8978 10652 8984
rect 9956 8492 10008 8498
rect 9956 8434 10008 8440
rect 9968 8362 9996 8434
rect 9956 8356 10008 8362
rect 9956 8298 10008 8304
rect 9968 7750 9996 8298
rect 9956 7744 10008 7750
rect 9956 7686 10008 7692
rect 10600 7744 10652 7750
rect 10600 7686 10652 7692
rect 9772 7540 9824 7546
rect 9772 7482 9824 7488
rect 9680 7404 9732 7410
rect 9680 7346 9732 7352
rect 9588 7336 9640 7342
rect 9588 7278 9640 7284
rect 9600 7002 9628 7278
rect 9128 6996 9180 7002
rect 9128 6938 9180 6944
rect 9588 6996 9640 7002
rect 9588 6938 9640 6944
rect 9692 6798 9720 7346
rect 9784 6798 9812 7482
rect 10612 7478 10640 7686
rect 10600 7472 10652 7478
rect 10600 7414 10652 7420
rect 10704 7410 10732 10474
rect 10888 8294 10916 11018
rect 11164 9994 11192 11494
rect 11428 11280 11480 11286
rect 11428 11222 11480 11228
rect 11440 10606 11468 11222
rect 11532 11150 11560 14962
rect 11716 13977 11744 14962
rect 11900 14482 11928 14962
rect 11992 14618 12020 17138
rect 12176 16590 12204 17682
rect 12256 17672 12308 17678
rect 12256 17614 12308 17620
rect 12268 16590 12296 17614
rect 12636 16658 12664 18022
rect 12728 17218 12756 18362
rect 12820 18154 12848 20198
rect 12900 19712 12952 19718
rect 12900 19654 12952 19660
rect 12912 18766 12940 19654
rect 12900 18760 12952 18766
rect 12900 18702 12952 18708
rect 12912 18306 12940 18702
rect 13004 18698 13032 20810
rect 13096 20602 13124 20878
rect 13084 20596 13136 20602
rect 13084 20538 13136 20544
rect 13084 20324 13136 20330
rect 13084 20266 13136 20272
rect 13096 19922 13124 20266
rect 13280 19990 13308 22442
rect 13372 22030 13400 22578
rect 13728 22568 13780 22574
rect 13728 22510 13780 22516
rect 13740 22030 13768 22510
rect 13360 22024 13412 22030
rect 13360 21966 13412 21972
rect 13728 22024 13780 22030
rect 13728 21966 13780 21972
rect 13544 21888 13596 21894
rect 13544 21830 13596 21836
rect 13360 20800 13412 20806
rect 13360 20742 13412 20748
rect 13372 20466 13400 20742
rect 13556 20466 13584 21830
rect 13634 21584 13690 21593
rect 14108 21554 14136 22646
rect 14292 22438 14320 23122
rect 14280 22432 14332 22438
rect 14280 22374 14332 22380
rect 14292 22098 14320 22374
rect 14280 22092 14332 22098
rect 14280 22034 14332 22040
rect 14464 22024 14516 22030
rect 14464 21966 14516 21972
rect 14280 21956 14332 21962
rect 14280 21898 14332 21904
rect 14292 21554 14320 21898
rect 14372 21888 14424 21894
rect 14372 21830 14424 21836
rect 13634 21519 13636 21528
rect 13688 21519 13690 21528
rect 14096 21548 14148 21554
rect 13636 21490 13688 21496
rect 14096 21490 14148 21496
rect 14280 21548 14332 21554
rect 14280 21490 14332 21496
rect 13728 21412 13780 21418
rect 13728 21354 13780 21360
rect 13636 21344 13688 21350
rect 13636 21286 13688 21292
rect 13360 20460 13412 20466
rect 13360 20402 13412 20408
rect 13452 20460 13504 20466
rect 13452 20402 13504 20408
rect 13544 20460 13596 20466
rect 13544 20402 13596 20408
rect 13464 20262 13492 20402
rect 13452 20256 13504 20262
rect 13452 20198 13504 20204
rect 13464 20097 13492 20198
rect 13450 20088 13506 20097
rect 13450 20023 13506 20032
rect 13268 19984 13320 19990
rect 13268 19926 13320 19932
rect 13084 19916 13136 19922
rect 13084 19858 13136 19864
rect 13280 19854 13308 19926
rect 13268 19848 13320 19854
rect 13268 19790 13320 19796
rect 13452 19848 13504 19854
rect 13452 19790 13504 19796
rect 13280 19174 13308 19790
rect 13464 19258 13492 19790
rect 13648 19666 13676 21286
rect 13740 19854 13768 21354
rect 14004 21140 14056 21146
rect 14004 21082 14056 21088
rect 13912 20800 13964 20806
rect 13912 20742 13964 20748
rect 13924 20466 13952 20742
rect 13912 20460 13964 20466
rect 13912 20402 13964 20408
rect 13924 20369 13952 20402
rect 13910 20360 13966 20369
rect 13910 20295 13966 20304
rect 13728 19848 13780 19854
rect 13912 19848 13964 19854
rect 13728 19790 13780 19796
rect 13832 19808 13912 19836
rect 13648 19638 13768 19666
rect 13636 19508 13688 19514
rect 13636 19450 13688 19456
rect 13372 19242 13492 19258
rect 13360 19236 13492 19242
rect 13412 19230 13492 19236
rect 13360 19178 13412 19184
rect 13176 19168 13228 19174
rect 13176 19110 13228 19116
rect 13268 19168 13320 19174
rect 13268 19110 13320 19116
rect 13084 18760 13136 18766
rect 13084 18702 13136 18708
rect 12992 18692 13044 18698
rect 12992 18634 13044 18640
rect 12912 18278 13032 18306
rect 13004 18222 13032 18278
rect 12992 18216 13044 18222
rect 12992 18158 13044 18164
rect 12808 18148 12860 18154
rect 12808 18090 12860 18096
rect 13096 17882 13124 18702
rect 13188 18426 13216 19110
rect 13268 18624 13320 18630
rect 13268 18566 13320 18572
rect 13360 18624 13412 18630
rect 13360 18566 13412 18572
rect 13176 18420 13228 18426
rect 13176 18362 13228 18368
rect 13280 18290 13308 18566
rect 13176 18284 13228 18290
rect 13176 18226 13228 18232
rect 13268 18284 13320 18290
rect 13268 18226 13320 18232
rect 13084 17876 13136 17882
rect 13084 17818 13136 17824
rect 12992 17740 13044 17746
rect 12992 17682 13044 17688
rect 12808 17264 12860 17270
rect 12728 17212 12808 17218
rect 12728 17206 12860 17212
rect 12728 17190 12848 17206
rect 12624 16652 12676 16658
rect 12624 16594 12676 16600
rect 12164 16584 12216 16590
rect 12164 16526 12216 16532
rect 12256 16584 12308 16590
rect 12256 16526 12308 16532
rect 12624 15020 12676 15026
rect 12624 14962 12676 14968
rect 12256 14884 12308 14890
rect 12256 14826 12308 14832
rect 11980 14612 12032 14618
rect 11980 14554 12032 14560
rect 11888 14476 11940 14482
rect 11888 14418 11940 14424
rect 11900 14006 11928 14418
rect 12268 14278 12296 14826
rect 12636 14618 12664 14962
rect 12624 14612 12676 14618
rect 12624 14554 12676 14560
rect 12728 14482 12756 17190
rect 12900 16992 12952 16998
rect 12900 16934 12952 16940
rect 12912 16590 12940 16934
rect 12900 16584 12952 16590
rect 12900 16526 12952 16532
rect 12808 16448 12860 16454
rect 12808 16390 12860 16396
rect 12820 16182 12848 16390
rect 13004 16182 13032 17682
rect 12808 16176 12860 16182
rect 12808 16118 12860 16124
rect 12992 16176 13044 16182
rect 12992 16118 13044 16124
rect 12808 15904 12860 15910
rect 12808 15846 12860 15852
rect 12820 15162 12848 15846
rect 12808 15156 12860 15162
rect 12808 15098 12860 15104
rect 13188 14958 13216 18226
rect 13268 17672 13320 17678
rect 13268 17614 13320 17620
rect 13280 16998 13308 17614
rect 13268 16992 13320 16998
rect 13268 16934 13320 16940
rect 13280 16590 13308 16934
rect 13372 16658 13400 18566
rect 13452 17672 13504 17678
rect 13452 17614 13504 17620
rect 13464 17082 13492 17614
rect 13648 17202 13676 19450
rect 13740 19378 13768 19638
rect 13728 19372 13780 19378
rect 13728 19314 13780 19320
rect 13832 19310 13860 19808
rect 13912 19790 13964 19796
rect 14016 19514 14044 21082
rect 14188 20936 14240 20942
rect 14186 20904 14188 20913
rect 14240 20904 14242 20913
rect 14186 20839 14242 20848
rect 14096 20528 14148 20534
rect 14094 20496 14096 20505
rect 14148 20496 14150 20505
rect 14094 20431 14150 20440
rect 14004 19508 14056 19514
rect 14004 19450 14056 19456
rect 14200 19446 14228 20839
rect 14188 19440 14240 19446
rect 14188 19382 14240 19388
rect 13820 19304 13872 19310
rect 13820 19246 13872 19252
rect 13832 18834 13860 19246
rect 13820 18828 13872 18834
rect 13820 18770 13872 18776
rect 13636 17196 13688 17202
rect 13636 17138 13688 17144
rect 13544 17128 13596 17134
rect 13464 17076 13544 17082
rect 13464 17070 13596 17076
rect 13464 17054 13584 17070
rect 13464 16794 13492 17054
rect 13648 16794 13676 17138
rect 13832 16998 13860 18770
rect 14200 17746 14228 19382
rect 14188 17740 14240 17746
rect 14188 17682 14240 17688
rect 13912 17128 13964 17134
rect 13912 17070 13964 17076
rect 13820 16992 13872 16998
rect 13820 16934 13872 16940
rect 13452 16788 13504 16794
rect 13452 16730 13504 16736
rect 13636 16788 13688 16794
rect 13636 16730 13688 16736
rect 13360 16652 13412 16658
rect 13360 16594 13412 16600
rect 13268 16584 13320 16590
rect 13268 16526 13320 16532
rect 13636 15020 13688 15026
rect 13636 14962 13688 14968
rect 13176 14952 13228 14958
rect 13176 14894 13228 14900
rect 13452 14884 13504 14890
rect 13452 14826 13504 14832
rect 12716 14476 12768 14482
rect 12716 14418 12768 14424
rect 12900 14340 12952 14346
rect 12900 14282 12952 14288
rect 12256 14272 12308 14278
rect 12256 14214 12308 14220
rect 11888 14000 11940 14006
rect 11702 13968 11758 13977
rect 11888 13942 11940 13948
rect 11702 13903 11758 13912
rect 12268 13394 12296 14214
rect 12912 13938 12940 14282
rect 12992 14272 13044 14278
rect 12992 14214 13044 14220
rect 12900 13932 12952 13938
rect 12900 13874 12952 13880
rect 12808 13728 12860 13734
rect 12808 13670 12860 13676
rect 12256 13388 12308 13394
rect 12256 13330 12308 13336
rect 12820 13326 12848 13670
rect 13004 13326 13032 14214
rect 13464 14006 13492 14826
rect 13542 14512 13598 14521
rect 13542 14447 13598 14456
rect 13556 14414 13584 14447
rect 13648 14414 13676 14962
rect 13544 14408 13596 14414
rect 13544 14350 13596 14356
rect 13636 14408 13688 14414
rect 13636 14350 13688 14356
rect 13452 14000 13504 14006
rect 13452 13942 13504 13948
rect 13084 13932 13136 13938
rect 13084 13874 13136 13880
rect 12348 13320 12400 13326
rect 12716 13320 12768 13326
rect 12400 13268 12572 13274
rect 12348 13262 12572 13268
rect 12716 13262 12768 13268
rect 12808 13320 12860 13326
rect 12808 13262 12860 13268
rect 12992 13320 13044 13326
rect 12992 13262 13044 13268
rect 11704 13252 11756 13258
rect 12360 13246 12572 13262
rect 11704 13194 11756 13200
rect 11612 11212 11664 11218
rect 11612 11154 11664 11160
rect 11520 11144 11572 11150
rect 11520 11086 11572 11092
rect 11520 10668 11572 10674
rect 11520 10610 11572 10616
rect 11428 10600 11480 10606
rect 11428 10542 11480 10548
rect 11152 9988 11204 9994
rect 11152 9930 11204 9936
rect 11164 9722 11192 9930
rect 11440 9926 11468 10542
rect 11532 9994 11560 10610
rect 11624 10062 11652 11154
rect 11612 10056 11664 10062
rect 11612 9998 11664 10004
rect 11520 9988 11572 9994
rect 11520 9930 11572 9936
rect 11428 9920 11480 9926
rect 11428 9862 11480 9868
rect 11152 9716 11204 9722
rect 11152 9658 11204 9664
rect 10876 8288 10928 8294
rect 10876 8230 10928 8236
rect 10888 7478 10916 8230
rect 10876 7472 10928 7478
rect 10876 7414 10928 7420
rect 11624 7410 11652 9998
rect 11716 9178 11744 13194
rect 12164 13184 12216 13190
rect 12164 13126 12216 13132
rect 12176 12434 12204 13126
rect 12176 12406 12388 12434
rect 12256 11756 12308 11762
rect 12256 11698 12308 11704
rect 12164 11348 12216 11354
rect 12164 11290 12216 11296
rect 11888 11212 11940 11218
rect 11808 11172 11888 11200
rect 11808 10674 11836 11172
rect 11888 11154 11940 11160
rect 11980 11144 12032 11150
rect 11978 11112 11980 11121
rect 12032 11112 12034 11121
rect 11978 11047 12034 11056
rect 11980 11008 12032 11014
rect 11980 10950 12032 10956
rect 11992 10674 12020 10950
rect 12176 10674 12204 11290
rect 11796 10668 11848 10674
rect 11796 10610 11848 10616
rect 11888 10668 11940 10674
rect 11888 10610 11940 10616
rect 11980 10668 12032 10674
rect 11980 10610 12032 10616
rect 12164 10668 12216 10674
rect 12164 10610 12216 10616
rect 11900 10266 11928 10610
rect 11888 10260 11940 10266
rect 11888 10202 11940 10208
rect 12176 10130 12204 10610
rect 12164 10124 12216 10130
rect 12164 10066 12216 10072
rect 12072 10056 12124 10062
rect 12072 9998 12124 10004
rect 11704 9172 11756 9178
rect 11704 9114 11756 9120
rect 12084 8974 12112 9998
rect 12176 9926 12204 10066
rect 12164 9920 12216 9926
rect 12164 9862 12216 9868
rect 12268 9674 12296 11698
rect 12360 11150 12388 12406
rect 12452 11898 12480 13246
rect 12544 13190 12572 13246
rect 12532 13184 12584 13190
rect 12532 13126 12584 13132
rect 12728 12986 12756 13262
rect 12716 12980 12768 12986
rect 12716 12922 12768 12928
rect 12728 12458 12756 12922
rect 12820 12646 12848 13262
rect 13004 12918 13032 13262
rect 12992 12912 13044 12918
rect 12992 12854 13044 12860
rect 12808 12640 12860 12646
rect 12808 12582 12860 12588
rect 12728 12430 12848 12458
rect 13096 12434 13124 13874
rect 13728 13796 13780 13802
rect 13728 13738 13780 13744
rect 13542 13696 13598 13705
rect 13542 13631 13598 13640
rect 13556 13326 13584 13631
rect 13544 13320 13596 13326
rect 13544 13262 13596 13268
rect 13360 13184 13412 13190
rect 13360 13126 13412 13132
rect 13268 12640 13320 12646
rect 13268 12582 13320 12588
rect 12532 12232 12584 12238
rect 12532 12174 12584 12180
rect 12624 12232 12676 12238
rect 12624 12174 12676 12180
rect 12440 11892 12492 11898
rect 12440 11834 12492 11840
rect 12544 11354 12572 12174
rect 12636 11898 12664 12174
rect 12716 12164 12768 12170
rect 12716 12106 12768 12112
rect 12624 11892 12676 11898
rect 12624 11834 12676 11840
rect 12624 11688 12676 11694
rect 12624 11630 12676 11636
rect 12532 11348 12584 11354
rect 12532 11290 12584 11296
rect 12348 11144 12400 11150
rect 12636 11098 12664 11630
rect 12728 11150 12756 12106
rect 12348 11086 12400 11092
rect 12360 11014 12388 11086
rect 12544 11070 12664 11098
rect 12716 11144 12768 11150
rect 12716 11086 12768 11092
rect 12820 11098 12848 12430
rect 12912 12406 13124 12434
rect 12912 12306 12940 12406
rect 12900 12300 12952 12306
rect 12900 12242 12952 12248
rect 12912 11286 12940 12242
rect 13176 12232 13228 12238
rect 13176 12174 13228 12180
rect 12990 11928 13046 11937
rect 13188 11898 13216 12174
rect 12990 11863 12992 11872
rect 13044 11863 13046 11872
rect 13176 11892 13228 11898
rect 12992 11834 13044 11840
rect 13176 11834 13228 11840
rect 13084 11756 13136 11762
rect 13004 11716 13084 11744
rect 12900 11280 12952 11286
rect 12900 11222 12952 11228
rect 12898 11112 12954 11121
rect 12820 11070 12898 11098
rect 12348 11008 12400 11014
rect 12348 10950 12400 10956
rect 12544 9674 12572 11070
rect 12898 11047 12954 11056
rect 12624 11008 12676 11014
rect 12624 10950 12676 10956
rect 12636 10674 12664 10950
rect 12624 10668 12676 10674
rect 12624 10610 12676 10616
rect 12808 10668 12860 10674
rect 12808 10610 12860 10616
rect 12624 10464 12676 10470
rect 12624 10406 12676 10412
rect 12636 10062 12664 10406
rect 12624 10056 12676 10062
rect 12624 9998 12676 10004
rect 12716 10056 12768 10062
rect 12716 9998 12768 10004
rect 12728 9926 12756 9998
rect 12624 9920 12676 9926
rect 12624 9862 12676 9868
rect 12716 9920 12768 9926
rect 12716 9862 12768 9868
rect 12176 9646 12296 9674
rect 12452 9646 12572 9674
rect 12176 9586 12204 9646
rect 12164 9580 12216 9586
rect 12164 9522 12216 9528
rect 12256 9580 12308 9586
rect 12452 9568 12480 9646
rect 12636 9586 12664 9862
rect 12624 9580 12676 9586
rect 12308 9540 12572 9568
rect 12256 9522 12308 9528
rect 12072 8968 12124 8974
rect 12072 8910 12124 8916
rect 11704 8832 11756 8838
rect 11704 8774 11756 8780
rect 11716 8634 11744 8774
rect 11704 8628 11756 8634
rect 11704 8570 11756 8576
rect 10692 7404 10744 7410
rect 10692 7346 10744 7352
rect 11612 7404 11664 7410
rect 11612 7346 11664 7352
rect 11716 7342 11744 8570
rect 12176 7857 12204 9522
rect 12256 9376 12308 9382
rect 12256 9318 12308 9324
rect 12348 9376 12400 9382
rect 12348 9318 12400 9324
rect 12268 8974 12296 9318
rect 12360 8974 12388 9318
rect 12256 8968 12308 8974
rect 12256 8910 12308 8916
rect 12348 8968 12400 8974
rect 12348 8910 12400 8916
rect 12440 8832 12492 8838
rect 12440 8774 12492 8780
rect 12162 7848 12218 7857
rect 12162 7783 12218 7792
rect 12348 7812 12400 7818
rect 12176 7698 12204 7783
rect 12452 7800 12480 8774
rect 12544 7970 12572 9540
rect 12624 9522 12676 9528
rect 12714 9480 12770 9489
rect 12714 9415 12716 9424
rect 12768 9415 12770 9424
rect 12716 9386 12768 9392
rect 12820 9178 12848 10610
rect 12912 10062 12940 11047
rect 13004 11014 13032 11716
rect 13084 11698 13136 11704
rect 13176 11756 13228 11762
rect 13176 11698 13228 11704
rect 13188 11558 13216 11698
rect 13176 11552 13228 11558
rect 13176 11494 13228 11500
rect 13176 11348 13228 11354
rect 13176 11290 13228 11296
rect 13084 11212 13136 11218
rect 13084 11154 13136 11160
rect 12992 11008 13044 11014
rect 12992 10950 13044 10956
rect 13004 10674 13032 10950
rect 12992 10668 13044 10674
rect 12992 10610 13044 10616
rect 13096 10266 13124 11154
rect 12992 10260 13044 10266
rect 12992 10202 13044 10208
rect 13084 10260 13136 10266
rect 13084 10202 13136 10208
rect 13004 10146 13032 10202
rect 13004 10118 13124 10146
rect 12900 10056 12952 10062
rect 12900 9998 12952 10004
rect 12912 9568 12940 9998
rect 12992 9580 13044 9586
rect 12912 9540 12992 9568
rect 12992 9522 13044 9528
rect 13096 9466 13124 10118
rect 12900 9444 12952 9450
rect 12900 9386 12952 9392
rect 13004 9438 13124 9466
rect 12808 9172 12860 9178
rect 12808 9114 12860 9120
rect 12624 9104 12676 9110
rect 12624 9046 12676 9052
rect 12636 8090 12664 9046
rect 12808 8492 12860 8498
rect 12808 8434 12860 8440
rect 12624 8084 12676 8090
rect 12624 8026 12676 8032
rect 12544 7942 12664 7970
rect 12532 7880 12584 7886
rect 12532 7822 12584 7828
rect 12400 7772 12480 7800
rect 12348 7754 12400 7760
rect 12176 7670 12296 7698
rect 12162 7576 12218 7585
rect 12162 7511 12164 7520
rect 12216 7511 12218 7520
rect 12164 7482 12216 7488
rect 11888 7404 11940 7410
rect 11888 7346 11940 7352
rect 11704 7336 11756 7342
rect 11704 7278 11756 7284
rect 11900 6934 11928 7346
rect 12268 6934 12296 7670
rect 12452 7478 12480 7772
rect 12440 7472 12492 7478
rect 12440 7414 12492 7420
rect 12440 7200 12492 7206
rect 12440 7142 12492 7148
rect 11888 6928 11940 6934
rect 11888 6870 11940 6876
rect 12256 6928 12308 6934
rect 12256 6870 12308 6876
rect 9680 6792 9732 6798
rect 9680 6734 9732 6740
rect 9772 6792 9824 6798
rect 9772 6734 9824 6740
rect 10324 6792 10376 6798
rect 10324 6734 10376 6740
rect 9692 6254 9720 6734
rect 10232 6656 10284 6662
rect 10232 6598 10284 6604
rect 10244 6322 10272 6598
rect 10232 6316 10284 6322
rect 10232 6258 10284 6264
rect 10336 6254 10364 6734
rect 11900 6390 11928 6870
rect 12452 6798 12480 7142
rect 12440 6792 12492 6798
rect 12440 6734 12492 6740
rect 12544 6458 12572 7822
rect 12636 7177 12664 7942
rect 12716 7880 12768 7886
rect 12716 7822 12768 7828
rect 12622 7168 12678 7177
rect 12622 7103 12678 7112
rect 12636 6934 12664 7103
rect 12624 6928 12676 6934
rect 12624 6870 12676 6876
rect 12728 6662 12756 7822
rect 12820 6882 12848 8434
rect 12912 8106 12940 9386
rect 13004 9110 13032 9438
rect 13188 9364 13216 11290
rect 13280 11150 13308 12582
rect 13372 11898 13400 13126
rect 13544 12844 13596 12850
rect 13544 12786 13596 12792
rect 13360 11892 13412 11898
rect 13360 11834 13412 11840
rect 13556 11558 13584 12786
rect 13740 12434 13768 13738
rect 13820 13728 13872 13734
rect 13820 13670 13872 13676
rect 13832 13530 13860 13670
rect 13820 13524 13872 13530
rect 13820 13466 13872 13472
rect 13924 13394 13952 17070
rect 14004 14952 14056 14958
rect 14004 14894 14056 14900
rect 14016 13394 14044 14894
rect 14200 14822 14228 17682
rect 14292 15026 14320 21490
rect 14384 21418 14412 21830
rect 14476 21690 14504 21966
rect 14464 21684 14516 21690
rect 14464 21626 14516 21632
rect 14372 21412 14424 21418
rect 14372 21354 14424 21360
rect 14384 20942 14412 21354
rect 14372 20936 14424 20942
rect 14372 20878 14424 20884
rect 14568 20466 14596 23666
rect 15384 23520 15436 23526
rect 15384 23462 15436 23468
rect 15200 21888 15252 21894
rect 15200 21830 15252 21836
rect 14924 21548 14976 21554
rect 14924 21490 14976 21496
rect 15108 21548 15160 21554
rect 15108 21490 15160 21496
rect 14648 20936 14700 20942
rect 14648 20878 14700 20884
rect 14556 20460 14608 20466
rect 14556 20402 14608 20408
rect 14372 20392 14424 20398
rect 14372 20334 14424 20340
rect 14384 19854 14412 20334
rect 14568 19854 14596 20402
rect 14660 19990 14688 20878
rect 14936 20058 14964 21490
rect 15120 21078 15148 21490
rect 15108 21072 15160 21078
rect 15028 21020 15108 21026
rect 15028 21014 15160 21020
rect 15028 20998 15148 21014
rect 15212 21010 15240 21830
rect 15200 21004 15252 21010
rect 15028 20602 15056 20998
rect 15200 20946 15252 20952
rect 15108 20936 15160 20942
rect 15108 20878 15160 20884
rect 15016 20596 15068 20602
rect 15016 20538 15068 20544
rect 14924 20052 14976 20058
rect 14924 19994 14976 20000
rect 14648 19984 14700 19990
rect 14648 19926 14700 19932
rect 15028 19922 15056 20538
rect 15016 19916 15068 19922
rect 15016 19858 15068 19864
rect 15120 19854 15148 20878
rect 15212 20058 15240 20946
rect 15396 20466 15424 23462
rect 15476 20868 15528 20874
rect 15476 20810 15528 20816
rect 15292 20460 15344 20466
rect 15292 20402 15344 20408
rect 15384 20460 15436 20466
rect 15384 20402 15436 20408
rect 15200 20052 15252 20058
rect 15200 19994 15252 20000
rect 14372 19848 14424 19854
rect 14372 19790 14424 19796
rect 14556 19848 14608 19854
rect 15108 19848 15160 19854
rect 14608 19808 14780 19836
rect 14556 19790 14608 19796
rect 14752 18766 14780 19808
rect 15108 19790 15160 19796
rect 15120 18970 15148 19790
rect 15200 19236 15252 19242
rect 15200 19178 15252 19184
rect 15108 18964 15160 18970
rect 15108 18906 15160 18912
rect 15108 18828 15160 18834
rect 15108 18770 15160 18776
rect 14648 18760 14700 18766
rect 14648 18702 14700 18708
rect 14740 18760 14792 18766
rect 14740 18702 14792 18708
rect 14660 18170 14688 18702
rect 14752 18306 14780 18702
rect 14752 18278 14872 18306
rect 14660 18142 14780 18170
rect 14752 18086 14780 18142
rect 14740 18080 14792 18086
rect 14740 18022 14792 18028
rect 14464 17536 14516 17542
rect 14464 17478 14516 17484
rect 14556 17536 14608 17542
rect 14556 17478 14608 17484
rect 14476 17270 14504 17478
rect 14464 17264 14516 17270
rect 14464 17206 14516 17212
rect 14568 17202 14596 17478
rect 14752 17202 14780 18022
rect 14844 17678 14872 18278
rect 15016 18080 15068 18086
rect 15016 18022 15068 18028
rect 15028 17814 15056 18022
rect 15016 17808 15068 17814
rect 15016 17750 15068 17756
rect 14832 17672 14884 17678
rect 14832 17614 14884 17620
rect 15016 17672 15068 17678
rect 15120 17660 15148 18770
rect 15212 18766 15240 19178
rect 15304 18970 15332 20402
rect 15292 18964 15344 18970
rect 15292 18906 15344 18912
rect 15200 18760 15252 18766
rect 15200 18702 15252 18708
rect 15304 18290 15332 18906
rect 15396 18358 15424 20402
rect 15488 20058 15516 20810
rect 15580 20602 15608 24074
rect 15764 23730 15792 24550
rect 15948 23730 15976 24550
rect 16212 24404 16264 24410
rect 16212 24346 16264 24352
rect 16224 24070 16252 24346
rect 16212 24064 16264 24070
rect 16212 24006 16264 24012
rect 15752 23724 15804 23730
rect 15752 23666 15804 23672
rect 15936 23724 15988 23730
rect 15936 23666 15988 23672
rect 16316 23526 16344 24754
rect 16592 24070 16620 24754
rect 17500 24744 17552 24750
rect 17500 24686 17552 24692
rect 17316 24608 17368 24614
rect 17316 24550 17368 24556
rect 17328 24342 17356 24550
rect 17316 24336 17368 24342
rect 17316 24278 17368 24284
rect 17224 24200 17276 24206
rect 16946 24168 17002 24177
rect 17224 24142 17276 24148
rect 16946 24103 16948 24112
rect 17000 24103 17002 24112
rect 16948 24074 17000 24080
rect 16488 24064 16540 24070
rect 16488 24006 16540 24012
rect 16580 24064 16632 24070
rect 16580 24006 16632 24012
rect 17132 24064 17184 24070
rect 17132 24006 17184 24012
rect 16396 23860 16448 23866
rect 16396 23802 16448 23808
rect 16408 23526 16436 23802
rect 16500 23526 16528 24006
rect 16592 23730 16620 24006
rect 16580 23724 16632 23730
rect 16580 23666 16632 23672
rect 15936 23520 15988 23526
rect 15936 23462 15988 23468
rect 16304 23520 16356 23526
rect 16304 23462 16356 23468
rect 16396 23520 16448 23526
rect 16396 23462 16448 23468
rect 16488 23520 16540 23526
rect 16488 23462 16540 23468
rect 15844 20800 15896 20806
rect 15844 20742 15896 20748
rect 15568 20596 15620 20602
rect 15568 20538 15620 20544
rect 15476 20052 15528 20058
rect 15476 19994 15528 20000
rect 15568 19508 15620 19514
rect 15568 19450 15620 19456
rect 15476 18896 15528 18902
rect 15476 18838 15528 18844
rect 15384 18352 15436 18358
rect 15384 18294 15436 18300
rect 15292 18284 15344 18290
rect 15292 18226 15344 18232
rect 15488 18222 15516 18838
rect 15476 18216 15528 18222
rect 15476 18158 15528 18164
rect 15068 17632 15148 17660
rect 15016 17614 15068 17620
rect 15028 17338 15056 17614
rect 15016 17332 15068 17338
rect 15016 17274 15068 17280
rect 14556 17196 14608 17202
rect 14556 17138 14608 17144
rect 14740 17196 14792 17202
rect 14740 17138 14792 17144
rect 14832 16992 14884 16998
rect 14832 16934 14884 16940
rect 15384 16992 15436 16998
rect 15384 16934 15436 16940
rect 14844 15162 14872 16934
rect 15396 16658 15424 16934
rect 15384 16652 15436 16658
rect 15384 16594 15436 16600
rect 15488 16522 15516 18158
rect 15476 16516 15528 16522
rect 15476 16458 15528 16464
rect 14832 15156 14884 15162
rect 14832 15098 14884 15104
rect 14280 15020 14332 15026
rect 14280 14962 14332 14968
rect 15200 14952 15252 14958
rect 15200 14894 15252 14900
rect 15292 14952 15344 14958
rect 15292 14894 15344 14900
rect 14188 14816 14240 14822
rect 14188 14758 14240 14764
rect 14200 14618 14228 14758
rect 14188 14612 14240 14618
rect 14188 14554 14240 14560
rect 15108 14612 15160 14618
rect 15108 14554 15160 14560
rect 14832 14408 14884 14414
rect 14832 14350 14884 14356
rect 15016 14408 15068 14414
rect 15016 14350 15068 14356
rect 14648 14272 14700 14278
rect 14648 14214 14700 14220
rect 14660 14006 14688 14214
rect 14648 14000 14700 14006
rect 14648 13942 14700 13948
rect 14096 13932 14148 13938
rect 14096 13874 14148 13880
rect 13912 13388 13964 13394
rect 13912 13330 13964 13336
rect 14004 13388 14056 13394
rect 14004 13330 14056 13336
rect 14108 13190 14136 13874
rect 14740 13728 14792 13734
rect 14740 13670 14792 13676
rect 14648 13320 14700 13326
rect 14752 13308 14780 13670
rect 14844 13530 14872 14350
rect 14832 13524 14884 13530
rect 14832 13466 14884 13472
rect 14924 13320 14976 13326
rect 14752 13280 14924 13308
rect 14648 13262 14700 13268
rect 14924 13262 14976 13268
rect 14096 13184 14148 13190
rect 14096 13126 14148 13132
rect 13648 12406 13768 12434
rect 13452 11552 13504 11558
rect 13452 11494 13504 11500
rect 13544 11552 13596 11558
rect 13544 11494 13596 11500
rect 13268 11144 13320 11150
rect 13268 11086 13320 11092
rect 13268 10600 13320 10606
rect 13268 10542 13320 10548
rect 13280 10266 13308 10542
rect 13464 10470 13492 11494
rect 13556 11150 13584 11494
rect 13648 11354 13676 12406
rect 13740 12374 13768 12406
rect 13728 12368 13780 12374
rect 13728 12310 13780 12316
rect 14108 12306 14136 13126
rect 14660 12850 14688 13262
rect 14936 12918 14964 13262
rect 14924 12912 14976 12918
rect 14924 12854 14976 12860
rect 14648 12844 14700 12850
rect 14648 12786 14700 12792
rect 14096 12300 14148 12306
rect 14096 12242 14148 12248
rect 14660 11898 14688 12786
rect 14648 11892 14700 11898
rect 14648 11834 14700 11840
rect 13912 11824 13964 11830
rect 13912 11766 13964 11772
rect 13820 11756 13872 11762
rect 13820 11698 13872 11704
rect 13728 11688 13780 11694
rect 13728 11630 13780 11636
rect 13636 11348 13688 11354
rect 13636 11290 13688 11296
rect 13636 11212 13688 11218
rect 13636 11154 13688 11160
rect 13544 11144 13596 11150
rect 13544 11086 13596 11092
rect 13452 10464 13504 10470
rect 13452 10406 13504 10412
rect 13268 10260 13320 10266
rect 13268 10202 13320 10208
rect 13544 10192 13596 10198
rect 13544 10134 13596 10140
rect 13556 10062 13584 10134
rect 13452 10056 13504 10062
rect 13452 9998 13504 10004
rect 13544 10056 13596 10062
rect 13544 9998 13596 10004
rect 13464 9586 13492 9998
rect 13556 9586 13584 9998
rect 13452 9580 13504 9586
rect 13372 9540 13452 9568
rect 13268 9376 13320 9382
rect 13188 9336 13268 9364
rect 13268 9318 13320 9324
rect 12992 9104 13044 9110
rect 12992 9046 13044 9052
rect 13084 8968 13136 8974
rect 13084 8910 13136 8916
rect 13096 8566 13124 8910
rect 13084 8560 13136 8566
rect 13084 8502 13136 8508
rect 13174 8120 13230 8129
rect 12912 8078 13124 8106
rect 12900 7880 12952 7886
rect 12900 7822 12952 7828
rect 12992 7880 13044 7886
rect 12992 7822 13044 7828
rect 12912 7002 12940 7822
rect 13004 7546 13032 7822
rect 12992 7540 13044 7546
rect 12992 7482 13044 7488
rect 13004 7206 13032 7482
rect 13096 7478 13124 8078
rect 13174 8055 13176 8064
rect 13228 8055 13230 8064
rect 13176 8026 13228 8032
rect 13176 7744 13228 7750
rect 13176 7686 13228 7692
rect 13084 7472 13136 7478
rect 13084 7414 13136 7420
rect 12992 7200 13044 7206
rect 12992 7142 13044 7148
rect 13084 7200 13136 7206
rect 13084 7142 13136 7148
rect 13096 7002 13124 7142
rect 12900 6996 12952 7002
rect 12900 6938 12952 6944
rect 13084 6996 13136 7002
rect 13084 6938 13136 6944
rect 12820 6854 13032 6882
rect 13004 6798 13032 6854
rect 12900 6792 12952 6798
rect 12898 6760 12900 6769
rect 12992 6792 13044 6798
rect 12952 6760 12954 6769
rect 12992 6734 13044 6740
rect 12898 6695 12954 6704
rect 12716 6656 12768 6662
rect 12716 6598 12768 6604
rect 12532 6452 12584 6458
rect 12532 6394 12584 6400
rect 13188 6390 13216 7686
rect 13280 7206 13308 9318
rect 13372 7750 13400 9540
rect 13452 9522 13504 9528
rect 13544 9580 13596 9586
rect 13544 9522 13596 9528
rect 13648 9450 13676 11154
rect 13740 11150 13768 11630
rect 13832 11558 13860 11698
rect 13820 11552 13872 11558
rect 13820 11494 13872 11500
rect 13728 11144 13780 11150
rect 13728 11086 13780 11092
rect 13924 9926 13952 11766
rect 14464 11552 14516 11558
rect 14464 11494 14516 11500
rect 14004 11076 14056 11082
rect 14004 11018 14056 11024
rect 14016 10674 14044 11018
rect 14476 10674 14504 11494
rect 14004 10668 14056 10674
rect 14004 10610 14056 10616
rect 14464 10668 14516 10674
rect 14464 10610 14516 10616
rect 14740 10668 14792 10674
rect 14740 10610 14792 10616
rect 14016 10130 14044 10610
rect 14096 10532 14148 10538
rect 14096 10474 14148 10480
rect 14108 10198 14136 10474
rect 14476 10470 14504 10610
rect 14464 10464 14516 10470
rect 14464 10406 14516 10412
rect 14752 10266 14780 10610
rect 14740 10260 14792 10266
rect 14740 10202 14792 10208
rect 14096 10192 14148 10198
rect 14096 10134 14148 10140
rect 14004 10124 14056 10130
rect 14004 10066 14056 10072
rect 14372 10056 14424 10062
rect 14372 9998 14424 10004
rect 14096 9988 14148 9994
rect 14096 9930 14148 9936
rect 13912 9920 13964 9926
rect 13912 9862 13964 9868
rect 13728 9648 13780 9654
rect 13728 9590 13780 9596
rect 13636 9444 13688 9450
rect 13636 9386 13688 9392
rect 13740 8362 13768 9590
rect 14108 8974 14136 9930
rect 14096 8968 14148 8974
rect 14096 8910 14148 8916
rect 13912 8492 13964 8498
rect 13912 8434 13964 8440
rect 13820 8424 13872 8430
rect 13820 8366 13872 8372
rect 13452 8356 13504 8362
rect 13452 8298 13504 8304
rect 13728 8356 13780 8362
rect 13728 8298 13780 8304
rect 13360 7744 13412 7750
rect 13360 7686 13412 7692
rect 13372 7410 13400 7686
rect 13464 7410 13492 8298
rect 13832 7886 13860 8366
rect 13924 8090 13952 8434
rect 13912 8084 13964 8090
rect 13912 8026 13964 8032
rect 13820 7880 13872 7886
rect 13820 7822 13872 7828
rect 13728 7812 13780 7818
rect 13728 7754 13780 7760
rect 13360 7404 13412 7410
rect 13360 7346 13412 7352
rect 13452 7404 13504 7410
rect 13452 7346 13504 7352
rect 13740 7342 13768 7754
rect 13832 7410 13860 7822
rect 13924 7410 13952 8026
rect 14108 7546 14136 8910
rect 14384 8634 14412 9998
rect 14372 8628 14424 8634
rect 14372 8570 14424 8576
rect 14924 8492 14976 8498
rect 14924 8434 14976 8440
rect 14936 8362 14964 8434
rect 14924 8356 14976 8362
rect 14924 8298 14976 8304
rect 14188 7812 14240 7818
rect 14188 7754 14240 7760
rect 14200 7721 14228 7754
rect 14556 7744 14608 7750
rect 14186 7712 14242 7721
rect 14556 7686 14608 7692
rect 14186 7647 14242 7656
rect 14096 7540 14148 7546
rect 14096 7482 14148 7488
rect 13820 7404 13872 7410
rect 13820 7346 13872 7352
rect 13912 7404 13964 7410
rect 13912 7346 13964 7352
rect 13728 7336 13780 7342
rect 13728 7278 13780 7284
rect 13268 7200 13320 7206
rect 13268 7142 13320 7148
rect 13280 7041 13308 7142
rect 13266 7032 13322 7041
rect 13266 6967 13322 6976
rect 13740 6798 13768 7278
rect 13268 6792 13320 6798
rect 13268 6734 13320 6740
rect 13728 6792 13780 6798
rect 13728 6734 13780 6740
rect 11888 6384 11940 6390
rect 11888 6326 11940 6332
rect 13176 6384 13228 6390
rect 13176 6326 13228 6332
rect 9680 6248 9732 6254
rect 9680 6190 9732 6196
rect 10324 6248 10376 6254
rect 10324 6190 10376 6196
rect 13280 5914 13308 6734
rect 13452 6724 13504 6730
rect 13452 6666 13504 6672
rect 13464 6322 13492 6666
rect 13740 6322 13768 6734
rect 13452 6316 13504 6322
rect 13452 6258 13504 6264
rect 13728 6316 13780 6322
rect 13728 6258 13780 6264
rect 13832 6186 13860 7346
rect 13924 7313 13952 7346
rect 13910 7304 13966 7313
rect 13910 7239 13966 7248
rect 14200 6866 14228 7647
rect 14568 7546 14596 7686
rect 14556 7540 14608 7546
rect 14556 7482 14608 7488
rect 14740 7472 14792 7478
rect 14660 7432 14740 7460
rect 14660 7426 14688 7432
rect 14568 7410 14688 7426
rect 14740 7414 14792 7420
rect 14830 7440 14886 7449
rect 14556 7404 14688 7410
rect 14608 7398 14688 7404
rect 14830 7375 14832 7384
rect 14556 7346 14608 7352
rect 14884 7375 14886 7384
rect 14832 7346 14884 7352
rect 14278 7304 14334 7313
rect 14278 7239 14334 7248
rect 14372 7268 14424 7274
rect 14188 6860 14240 6866
rect 14188 6802 14240 6808
rect 14292 6798 14320 7239
rect 14372 7210 14424 7216
rect 14384 6934 14412 7210
rect 14372 6928 14424 6934
rect 14372 6870 14424 6876
rect 14936 6798 14964 8298
rect 15028 7546 15056 14350
rect 15120 13326 15148 14554
rect 15108 13320 15160 13326
rect 15108 13262 15160 13268
rect 15212 12434 15240 14894
rect 15304 14498 15332 14894
rect 15488 14634 15516 16458
rect 15580 14822 15608 19450
rect 15856 19417 15884 20742
rect 15842 19408 15898 19417
rect 15842 19343 15898 19352
rect 15752 18760 15804 18766
rect 15752 18702 15804 18708
rect 15844 18760 15896 18766
rect 15844 18702 15896 18708
rect 15660 18148 15712 18154
rect 15660 18090 15712 18096
rect 15672 17762 15700 18090
rect 15764 17882 15792 18702
rect 15856 18290 15884 18702
rect 15844 18284 15896 18290
rect 15844 18226 15896 18232
rect 15752 17876 15804 17882
rect 15752 17818 15804 17824
rect 15672 17734 15792 17762
rect 15660 16992 15712 16998
rect 15660 16934 15712 16940
rect 15568 14816 15620 14822
rect 15568 14758 15620 14764
rect 15488 14606 15608 14634
rect 15672 14618 15700 16934
rect 15764 16574 15792 17734
rect 15842 17232 15898 17241
rect 15842 17167 15844 17176
rect 15896 17167 15898 17176
rect 15844 17138 15896 17144
rect 15856 16726 15884 17138
rect 15948 17105 15976 23462
rect 16120 22432 16172 22438
rect 16120 22374 16172 22380
rect 16132 21894 16160 22374
rect 16212 22160 16264 22166
rect 16212 22102 16264 22108
rect 16120 21888 16172 21894
rect 16120 21830 16172 21836
rect 16132 21554 16160 21830
rect 16120 21548 16172 21554
rect 16120 21490 16172 21496
rect 16028 21344 16080 21350
rect 16028 21286 16080 21292
rect 16040 19360 16068 21286
rect 16132 20942 16160 21490
rect 16224 21486 16252 22102
rect 16304 21956 16356 21962
rect 16304 21898 16356 21904
rect 16316 21554 16344 21898
rect 16304 21548 16356 21554
rect 16304 21490 16356 21496
rect 16212 21480 16264 21486
rect 16212 21422 16264 21428
rect 16224 21010 16252 21422
rect 16316 21146 16344 21490
rect 16304 21140 16356 21146
rect 16304 21082 16356 21088
rect 16212 21004 16264 21010
rect 16212 20946 16264 20952
rect 16120 20936 16172 20942
rect 16120 20878 16172 20884
rect 16316 20534 16344 21082
rect 16408 20602 16436 23462
rect 16592 22710 16620 23666
rect 16580 22704 16632 22710
rect 16580 22646 16632 22652
rect 17040 22094 17092 22098
rect 17144 22094 17172 24006
rect 17236 23662 17264 24142
rect 17328 23866 17356 24278
rect 17512 24188 17540 24686
rect 17776 24608 17828 24614
rect 17776 24550 17828 24556
rect 17788 24206 17816 24550
rect 18144 24404 18196 24410
rect 18144 24346 18196 24352
rect 18604 24404 18656 24410
rect 18604 24346 18656 24352
rect 17960 24336 18012 24342
rect 17960 24278 18012 24284
rect 17592 24200 17644 24206
rect 17512 24160 17592 24188
rect 17316 23860 17368 23866
rect 17316 23802 17368 23808
rect 17408 23792 17460 23798
rect 17408 23734 17460 23740
rect 17224 23656 17276 23662
rect 17224 23598 17276 23604
rect 17420 23610 17448 23734
rect 17512 23730 17540 24160
rect 17592 24142 17644 24148
rect 17684 24200 17736 24206
rect 17684 24142 17736 24148
rect 17776 24200 17828 24206
rect 17776 24142 17828 24148
rect 17500 23724 17552 23730
rect 17500 23666 17552 23672
rect 17420 23582 17632 23610
rect 17696 23594 17724 24142
rect 17868 24064 17920 24070
rect 17868 24006 17920 24012
rect 17880 23866 17908 24006
rect 17868 23860 17920 23866
rect 17868 23802 17920 23808
rect 17868 23724 17920 23730
rect 17868 23666 17920 23672
rect 17604 23526 17632 23582
rect 17684 23588 17736 23594
rect 17684 23530 17736 23536
rect 17500 23520 17552 23526
rect 17500 23462 17552 23468
rect 17592 23520 17644 23526
rect 17592 23462 17644 23468
rect 17316 22772 17368 22778
rect 17316 22714 17368 22720
rect 17224 22432 17276 22438
rect 17224 22374 17276 22380
rect 17040 22092 17172 22094
rect 17092 22066 17172 22092
rect 17040 22034 17092 22040
rect 17236 22030 17264 22374
rect 17328 22030 17356 22714
rect 17224 22024 17276 22030
rect 17224 21966 17276 21972
rect 17316 22024 17368 22030
rect 17316 21966 17368 21972
rect 17132 21888 17184 21894
rect 17132 21830 17184 21836
rect 17144 21554 17172 21830
rect 17328 21593 17356 21966
rect 17314 21584 17370 21593
rect 17132 21548 17184 21554
rect 17314 21519 17370 21528
rect 17132 21490 17184 21496
rect 17144 21010 17172 21490
rect 17408 21480 17460 21486
rect 17408 21422 17460 21428
rect 17224 21412 17276 21418
rect 17224 21354 17276 21360
rect 17132 21004 17184 21010
rect 17132 20946 17184 20952
rect 16580 20936 16632 20942
rect 16580 20878 16632 20884
rect 16396 20596 16448 20602
rect 16396 20538 16448 20544
rect 16304 20528 16356 20534
rect 16304 20470 16356 20476
rect 16212 20460 16264 20466
rect 16212 20402 16264 20408
rect 16224 20058 16252 20402
rect 16212 20052 16264 20058
rect 16264 20012 16344 20040
rect 16212 19994 16264 20000
rect 16120 19372 16172 19378
rect 16040 19332 16120 19360
rect 16120 19314 16172 19320
rect 16028 18624 16080 18630
rect 16028 18566 16080 18572
rect 16040 18154 16068 18566
rect 16028 18148 16080 18154
rect 16028 18090 16080 18096
rect 16040 17746 16068 18090
rect 16028 17740 16080 17746
rect 16028 17682 16080 17688
rect 16028 17536 16080 17542
rect 16028 17478 16080 17484
rect 16040 17202 16068 17478
rect 16028 17196 16080 17202
rect 16028 17138 16080 17144
rect 15934 17096 15990 17105
rect 15934 17031 15990 17040
rect 15844 16720 15896 16726
rect 15844 16662 15896 16668
rect 15764 16546 15884 16574
rect 15304 14470 15516 14498
rect 15292 14408 15344 14414
rect 15292 14350 15344 14356
rect 15304 13530 15332 14350
rect 15384 13728 15436 13734
rect 15384 13670 15436 13676
rect 15292 13524 15344 13530
rect 15292 13466 15344 13472
rect 15292 13320 15344 13326
rect 15292 13262 15344 13268
rect 15304 12646 15332 13262
rect 15396 12850 15424 13670
rect 15384 12844 15436 12850
rect 15384 12786 15436 12792
rect 15292 12640 15344 12646
rect 15292 12582 15344 12588
rect 15396 12442 15424 12786
rect 15384 12436 15436 12442
rect 15212 12406 15332 12434
rect 15200 11552 15252 11558
rect 15200 11494 15252 11500
rect 15212 11218 15240 11494
rect 15200 11212 15252 11218
rect 15200 11154 15252 11160
rect 15304 8129 15332 12406
rect 15384 12378 15436 12384
rect 15384 12164 15436 12170
rect 15384 12106 15436 12112
rect 15396 11150 15424 12106
rect 15488 11898 15516 14470
rect 15580 13530 15608 14606
rect 15660 14612 15712 14618
rect 15660 14554 15712 14560
rect 15660 14408 15712 14414
rect 15660 14350 15712 14356
rect 15672 14278 15700 14350
rect 15660 14272 15712 14278
rect 15660 14214 15712 14220
rect 15672 13818 15700 14214
rect 15856 13818 15884 16546
rect 16028 16448 16080 16454
rect 16028 16390 16080 16396
rect 15936 14816 15988 14822
rect 15936 14758 15988 14764
rect 15948 13938 15976 14758
rect 15936 13932 15988 13938
rect 15936 13874 15988 13880
rect 15934 13832 15990 13841
rect 15672 13790 15792 13818
rect 15856 13790 15934 13818
rect 15568 13524 15620 13530
rect 15568 13466 15620 13472
rect 15660 13320 15712 13326
rect 15660 13262 15712 13268
rect 15568 12844 15620 12850
rect 15568 12786 15620 12792
rect 15580 12170 15608 12786
rect 15672 12646 15700 13262
rect 15660 12640 15712 12646
rect 15660 12582 15712 12588
rect 15568 12164 15620 12170
rect 15568 12106 15620 12112
rect 15566 11928 15622 11937
rect 15476 11892 15528 11898
rect 15566 11863 15568 11872
rect 15476 11834 15528 11840
rect 15620 11863 15622 11872
rect 15568 11834 15620 11840
rect 15568 11756 15620 11762
rect 15568 11698 15620 11704
rect 15476 11688 15528 11694
rect 15476 11630 15528 11636
rect 15488 11286 15516 11630
rect 15476 11280 15528 11286
rect 15476 11222 15528 11228
rect 15384 11144 15436 11150
rect 15580 11121 15608 11698
rect 15672 11150 15700 12582
rect 15764 11150 15792 13790
rect 15934 13767 15990 13776
rect 15844 13524 15896 13530
rect 15844 13466 15896 13472
rect 15856 13394 15884 13466
rect 15948 13394 15976 13767
rect 15844 13388 15896 13394
rect 15844 13330 15896 13336
rect 15936 13388 15988 13394
rect 15936 13330 15988 13336
rect 16040 13190 16068 16390
rect 16028 13184 16080 13190
rect 16028 13126 16080 13132
rect 15842 13016 15898 13025
rect 15842 12951 15898 12960
rect 15856 12918 15884 12951
rect 15844 12912 15896 12918
rect 15844 12854 15896 12860
rect 16132 12850 16160 19314
rect 16316 17746 16344 20012
rect 16408 19854 16436 20538
rect 16396 19848 16448 19854
rect 16396 19790 16448 19796
rect 16592 19786 16620 20878
rect 17040 20460 17092 20466
rect 17040 20402 17092 20408
rect 16580 19780 16632 19786
rect 16580 19722 16632 19728
rect 16764 19780 16816 19786
rect 16764 19722 16816 19728
rect 16396 19712 16448 19718
rect 16396 19654 16448 19660
rect 16408 19446 16436 19654
rect 16396 19440 16448 19446
rect 16396 19382 16448 19388
rect 16408 18290 16436 19382
rect 16396 18284 16448 18290
rect 16396 18226 16448 18232
rect 16488 18080 16540 18086
rect 16488 18022 16540 18028
rect 16304 17740 16356 17746
rect 16304 17682 16356 17688
rect 16316 17202 16344 17682
rect 16396 17672 16448 17678
rect 16396 17614 16448 17620
rect 16212 17196 16264 17202
rect 16212 17138 16264 17144
rect 16304 17196 16356 17202
rect 16304 17138 16356 17144
rect 16224 17105 16252 17138
rect 16210 17096 16266 17105
rect 16210 17031 16266 17040
rect 16408 16726 16436 17614
rect 16500 16998 16528 18022
rect 16672 17808 16724 17814
rect 16672 17750 16724 17756
rect 16580 17604 16632 17610
rect 16580 17546 16632 17552
rect 16592 17338 16620 17546
rect 16684 17542 16712 17750
rect 16672 17536 16724 17542
rect 16672 17478 16724 17484
rect 16580 17332 16632 17338
rect 16580 17274 16632 17280
rect 16672 17196 16724 17202
rect 16672 17138 16724 17144
rect 16488 16992 16540 16998
rect 16488 16934 16540 16940
rect 16396 16720 16448 16726
rect 16684 16697 16712 17138
rect 16396 16662 16448 16668
rect 16670 16688 16726 16697
rect 16670 16623 16726 16632
rect 16684 16250 16712 16623
rect 16672 16244 16724 16250
rect 16672 16186 16724 16192
rect 16776 15858 16804 19722
rect 17052 18902 17080 20402
rect 17132 20324 17184 20330
rect 17132 20266 17184 20272
rect 17040 18896 17092 18902
rect 17040 18838 17092 18844
rect 17144 17678 17172 20266
rect 17236 19786 17264 21354
rect 17420 21010 17448 21422
rect 17408 21004 17460 21010
rect 17408 20946 17460 20952
rect 17314 20360 17370 20369
rect 17314 20295 17316 20304
rect 17368 20295 17370 20304
rect 17316 20266 17368 20272
rect 17224 19780 17276 19786
rect 17224 19722 17276 19728
rect 16948 17672 17000 17678
rect 16946 17640 16948 17649
rect 17132 17672 17184 17678
rect 17000 17640 17002 17649
rect 17132 17614 17184 17620
rect 16946 17575 17002 17584
rect 17224 17604 17276 17610
rect 17224 17546 17276 17552
rect 17316 17604 17368 17610
rect 17316 17546 17368 17552
rect 16856 17536 16908 17542
rect 16856 17478 16908 17484
rect 16868 16046 16896 17478
rect 16948 17196 17000 17202
rect 16948 17138 17000 17144
rect 17132 17196 17184 17202
rect 17132 17138 17184 17144
rect 16960 16250 16988 17138
rect 17040 17128 17092 17134
rect 17040 17070 17092 17076
rect 16948 16244 17000 16250
rect 16948 16186 17000 16192
rect 16856 16040 16908 16046
rect 16856 15982 16908 15988
rect 17052 15978 17080 17070
rect 17040 15972 17092 15978
rect 17040 15914 17092 15920
rect 16776 15830 16988 15858
rect 16960 15706 16988 15830
rect 16948 15700 17000 15706
rect 16948 15642 17000 15648
rect 16856 14952 16908 14958
rect 16856 14894 16908 14900
rect 16672 14408 16724 14414
rect 16672 14350 16724 14356
rect 16764 14408 16816 14414
rect 16764 14350 16816 14356
rect 16488 14068 16540 14074
rect 16488 14010 16540 14016
rect 16396 13252 16448 13258
rect 16396 13194 16448 13200
rect 16408 12986 16436 13194
rect 16396 12980 16448 12986
rect 16396 12922 16448 12928
rect 16120 12844 16172 12850
rect 16120 12786 16172 12792
rect 15844 12708 15896 12714
rect 15844 12650 15896 12656
rect 15856 12442 15884 12650
rect 15844 12436 15896 12442
rect 15844 12378 15896 12384
rect 15936 12436 15988 12442
rect 16408 12434 16436 12922
rect 15936 12378 15988 12384
rect 16224 12406 16436 12434
rect 15948 12322 15976 12378
rect 15856 12306 15976 12322
rect 15844 12300 15976 12306
rect 15896 12294 15976 12300
rect 15844 12242 15896 12248
rect 15844 12164 15896 12170
rect 15844 12106 15896 12112
rect 15856 11354 15884 12106
rect 15936 12096 15988 12102
rect 15936 12038 15988 12044
rect 15948 11762 15976 12038
rect 15936 11756 15988 11762
rect 15936 11698 15988 11704
rect 16120 11756 16172 11762
rect 16120 11698 16172 11704
rect 16132 11642 16160 11698
rect 15948 11614 16160 11642
rect 15844 11348 15896 11354
rect 15844 11290 15896 11296
rect 15948 11286 15976 11614
rect 16028 11552 16080 11558
rect 16028 11494 16080 11500
rect 15936 11280 15988 11286
rect 15936 11222 15988 11228
rect 16040 11150 16068 11494
rect 16224 11150 16252 12406
rect 16500 12238 16528 14010
rect 16580 14000 16632 14006
rect 16580 13942 16632 13948
rect 16592 12374 16620 13942
rect 16580 12368 16632 12374
rect 16580 12310 16632 12316
rect 16488 12232 16540 12238
rect 16488 12174 16540 12180
rect 16500 11762 16528 12174
rect 16580 12164 16632 12170
rect 16580 12106 16632 12112
rect 16304 11756 16356 11762
rect 16304 11698 16356 11704
rect 16488 11756 16540 11762
rect 16488 11698 16540 11704
rect 15660 11144 15712 11150
rect 15384 11086 15436 11092
rect 15566 11112 15622 11121
rect 15660 11086 15712 11092
rect 15752 11144 15804 11150
rect 16028 11144 16080 11150
rect 15752 11086 15804 11092
rect 15934 11112 15990 11121
rect 15566 11047 15622 11056
rect 16028 11086 16080 11092
rect 16212 11144 16264 11150
rect 16316 11121 16344 11698
rect 16396 11348 16448 11354
rect 16396 11290 16448 11296
rect 16212 11086 16264 11092
rect 16302 11112 16358 11121
rect 15934 11047 15990 11056
rect 15476 10804 15528 10810
rect 15476 10746 15528 10752
rect 15488 10713 15516 10746
rect 15948 10742 15976 11047
rect 15936 10736 15988 10742
rect 15474 10704 15530 10713
rect 15936 10678 15988 10684
rect 15474 10639 15530 10648
rect 15476 10600 15528 10606
rect 15476 10542 15528 10548
rect 15488 9994 15516 10542
rect 16040 10470 16068 11086
rect 16120 11008 16172 11014
rect 16120 10950 16172 10956
rect 16132 10674 16160 10950
rect 16120 10668 16172 10674
rect 16120 10610 16172 10616
rect 16028 10464 16080 10470
rect 16028 10406 16080 10412
rect 15476 9988 15528 9994
rect 15476 9930 15528 9936
rect 15290 8120 15346 8129
rect 15290 8055 15346 8064
rect 15200 7744 15252 7750
rect 15200 7686 15252 7692
rect 15016 7540 15068 7546
rect 15016 7482 15068 7488
rect 15212 7478 15240 7686
rect 15200 7472 15252 7478
rect 15200 7414 15252 7420
rect 15382 7440 15438 7449
rect 15108 7404 15160 7410
rect 15382 7375 15384 7384
rect 15108 7346 15160 7352
rect 15436 7375 15438 7384
rect 15384 7346 15436 7352
rect 15014 7032 15070 7041
rect 15120 7002 15148 7346
rect 15396 7002 15424 7346
rect 15014 6967 15016 6976
rect 15068 6967 15070 6976
rect 15108 6996 15160 7002
rect 15016 6938 15068 6944
rect 15108 6938 15160 6944
rect 15384 6996 15436 7002
rect 15384 6938 15436 6944
rect 15488 6798 15516 9930
rect 16224 8974 16252 11086
rect 16302 11047 16358 11056
rect 16408 10962 16436 11290
rect 16500 11082 16528 11698
rect 16488 11076 16540 11082
rect 16488 11018 16540 11024
rect 16316 10934 16436 10962
rect 16316 10810 16344 10934
rect 16304 10804 16356 10810
rect 16304 10746 16356 10752
rect 16304 10668 16356 10674
rect 16304 10610 16356 10616
rect 16316 9926 16344 10610
rect 16396 10464 16448 10470
rect 16396 10406 16448 10412
rect 16408 10266 16436 10406
rect 16396 10260 16448 10266
rect 16396 10202 16448 10208
rect 16304 9920 16356 9926
rect 16304 9862 16356 9868
rect 16212 8968 16264 8974
rect 16212 8910 16264 8916
rect 15936 8288 15988 8294
rect 15936 8230 15988 8236
rect 16120 8288 16172 8294
rect 16120 8230 16172 8236
rect 15948 7886 15976 8230
rect 16028 8016 16080 8022
rect 16028 7958 16080 7964
rect 15752 7880 15804 7886
rect 15936 7880 15988 7886
rect 15752 7822 15804 7828
rect 15842 7848 15898 7857
rect 15568 7404 15620 7410
rect 15568 7346 15620 7352
rect 15580 6934 15608 7346
rect 15764 7002 15792 7822
rect 15936 7822 15988 7828
rect 15842 7783 15898 7792
rect 15856 7410 15884 7783
rect 15948 7750 15976 7822
rect 15936 7744 15988 7750
rect 15936 7686 15988 7692
rect 15844 7404 15896 7410
rect 15844 7346 15896 7352
rect 15936 7404 15988 7410
rect 15936 7346 15988 7352
rect 15948 7177 15976 7346
rect 16040 7206 16068 7958
rect 16028 7200 16080 7206
rect 15934 7168 15990 7177
rect 16028 7142 16080 7148
rect 15934 7103 15990 7112
rect 15752 6996 15804 7002
rect 15752 6938 15804 6944
rect 15568 6928 15620 6934
rect 15568 6870 15620 6876
rect 15844 6928 15896 6934
rect 15844 6870 15896 6876
rect 15856 6798 15884 6870
rect 14280 6792 14332 6798
rect 14280 6734 14332 6740
rect 14924 6792 14976 6798
rect 14924 6734 14976 6740
rect 15476 6792 15528 6798
rect 15476 6734 15528 6740
rect 15844 6792 15896 6798
rect 15844 6734 15896 6740
rect 14292 6254 14320 6734
rect 14280 6248 14332 6254
rect 14280 6190 14332 6196
rect 13820 6180 13872 6186
rect 13820 6122 13872 6128
rect 15488 5914 15516 6734
rect 16040 6390 16068 7142
rect 16132 7041 16160 8230
rect 16210 7848 16266 7857
rect 16210 7783 16266 7792
rect 16224 7546 16252 7783
rect 16212 7540 16264 7546
rect 16212 7482 16264 7488
rect 16212 7404 16264 7410
rect 16212 7346 16264 7352
rect 16118 7032 16174 7041
rect 16118 6967 16174 6976
rect 16224 6730 16252 7346
rect 16316 7206 16344 9862
rect 16304 7200 16356 7206
rect 16304 7142 16356 7148
rect 16212 6724 16264 6730
rect 16212 6666 16264 6672
rect 16316 6662 16344 7142
rect 16500 6798 16528 11018
rect 16592 11014 16620 12106
rect 16580 11008 16632 11014
rect 16580 10950 16632 10956
rect 16684 10962 16712 14350
rect 16776 11937 16804 14350
rect 16868 13938 16896 14894
rect 16856 13932 16908 13938
rect 16856 13874 16908 13880
rect 16856 12300 16908 12306
rect 16856 12242 16908 12248
rect 16762 11928 16818 11937
rect 16762 11863 16818 11872
rect 16776 11558 16804 11863
rect 16764 11552 16816 11558
rect 16764 11494 16816 11500
rect 16592 10062 16620 10950
rect 16684 10934 16804 10962
rect 16672 10668 16724 10674
rect 16672 10610 16724 10616
rect 16684 10266 16712 10610
rect 16672 10260 16724 10266
rect 16672 10202 16724 10208
rect 16776 10198 16804 10934
rect 16764 10192 16816 10198
rect 16764 10134 16816 10140
rect 16580 10056 16632 10062
rect 16580 9998 16632 10004
rect 16592 9178 16620 9998
rect 16580 9172 16632 9178
rect 16580 9114 16632 9120
rect 16592 9042 16620 9114
rect 16580 9036 16632 9042
rect 16580 8978 16632 8984
rect 16868 8498 16896 12242
rect 16960 12170 16988 15642
rect 17144 14618 17172 17138
rect 17236 17105 17264 17546
rect 17328 17338 17356 17546
rect 17316 17332 17368 17338
rect 17316 17274 17368 17280
rect 17316 17128 17368 17134
rect 17222 17096 17278 17105
rect 17316 17070 17368 17076
rect 17222 17031 17278 17040
rect 17328 16726 17356 17070
rect 17512 16946 17540 23462
rect 17880 22778 17908 23666
rect 17972 23526 18000 24278
rect 18156 24274 18184 24346
rect 18144 24268 18196 24274
rect 18144 24210 18196 24216
rect 18616 24206 18644 24346
rect 19064 24268 19116 24274
rect 19064 24210 19116 24216
rect 19248 24268 19300 24274
rect 19248 24210 19300 24216
rect 18604 24200 18656 24206
rect 18050 24168 18106 24177
rect 18604 24142 18656 24148
rect 18050 24103 18106 24112
rect 18064 24070 18092 24103
rect 18052 24064 18104 24070
rect 18052 24006 18104 24012
rect 18616 23730 18644 24142
rect 18972 24132 19024 24138
rect 18972 24074 19024 24080
rect 18984 23866 19012 24074
rect 18972 23860 19024 23866
rect 18972 23802 19024 23808
rect 18604 23724 18656 23730
rect 18604 23666 18656 23672
rect 18880 23724 18932 23730
rect 18880 23666 18932 23672
rect 18512 23588 18564 23594
rect 18512 23530 18564 23536
rect 17960 23520 18012 23526
rect 17960 23462 18012 23468
rect 18052 23520 18104 23526
rect 18052 23462 18104 23468
rect 17868 22772 17920 22778
rect 17868 22714 17920 22720
rect 17684 21888 17736 21894
rect 17684 21830 17736 21836
rect 17696 20466 17724 21830
rect 17880 21486 17908 22714
rect 18064 21554 18092 23462
rect 18052 21548 18104 21554
rect 18052 21490 18104 21496
rect 17868 21480 17920 21486
rect 17868 21422 17920 21428
rect 17776 21412 17828 21418
rect 17776 21354 17828 21360
rect 17788 21010 17816 21354
rect 17880 21078 17908 21422
rect 17868 21072 17920 21078
rect 17868 21014 17920 21020
rect 17776 21004 17828 21010
rect 17776 20946 17828 20952
rect 17960 21004 18012 21010
rect 17960 20946 18012 20952
rect 17684 20460 17736 20466
rect 17684 20402 17736 20408
rect 17972 19922 18000 20946
rect 18064 20806 18092 21490
rect 18524 20874 18552 23530
rect 18616 22642 18644 23666
rect 18696 22976 18748 22982
rect 18696 22918 18748 22924
rect 18604 22636 18656 22642
rect 18604 22578 18656 22584
rect 18708 22094 18736 22918
rect 18708 22066 18828 22094
rect 18604 21072 18656 21078
rect 18604 21014 18656 21020
rect 18616 20942 18644 21014
rect 18604 20936 18656 20942
rect 18604 20878 18656 20884
rect 18328 20868 18380 20874
rect 18328 20810 18380 20816
rect 18512 20868 18564 20874
rect 18512 20810 18564 20816
rect 18052 20800 18104 20806
rect 18052 20742 18104 20748
rect 18236 20392 18288 20398
rect 18236 20334 18288 20340
rect 18248 20262 18276 20334
rect 18236 20256 18288 20262
rect 18236 20198 18288 20204
rect 18248 20058 18276 20198
rect 18236 20052 18288 20058
rect 18236 19994 18288 20000
rect 17960 19916 18012 19922
rect 17960 19858 18012 19864
rect 18144 19712 18196 19718
rect 18144 19654 18196 19660
rect 17776 18828 17828 18834
rect 17776 18770 17828 18776
rect 17788 18290 17816 18770
rect 17776 18284 17828 18290
rect 17696 18244 17776 18272
rect 17696 17202 17724 18244
rect 17776 18226 17828 18232
rect 17776 17672 17828 17678
rect 17776 17614 17828 17620
rect 17684 17196 17736 17202
rect 17684 17138 17736 17144
rect 17420 16918 17540 16946
rect 17316 16720 17368 16726
rect 17316 16662 17368 16668
rect 17224 16448 17276 16454
rect 17224 16390 17276 16396
rect 17132 14612 17184 14618
rect 17132 14554 17184 14560
rect 17236 14482 17264 16390
rect 17420 15978 17448 16918
rect 17500 16788 17552 16794
rect 17788 16776 17816 17614
rect 17868 17536 17920 17542
rect 17868 17478 17920 17484
rect 17960 17536 18012 17542
rect 17960 17478 18012 17484
rect 17880 16794 17908 17478
rect 17972 17270 18000 17478
rect 17960 17264 18012 17270
rect 17960 17206 18012 17212
rect 17552 16748 17816 16776
rect 17500 16730 17552 16736
rect 17788 16658 17816 16748
rect 17868 16788 17920 16794
rect 17868 16730 17920 16736
rect 17776 16652 17828 16658
rect 17776 16594 17828 16600
rect 18052 16584 18104 16590
rect 18050 16552 18052 16561
rect 18104 16552 18106 16561
rect 18050 16487 18106 16496
rect 18052 16448 18104 16454
rect 18052 16390 18104 16396
rect 18064 16114 18092 16390
rect 18052 16108 18104 16114
rect 18052 16050 18104 16056
rect 17960 16040 18012 16046
rect 17960 15982 18012 15988
rect 17408 15972 17460 15978
rect 17408 15914 17460 15920
rect 17040 14476 17092 14482
rect 17040 14418 17092 14424
rect 17224 14476 17276 14482
rect 17224 14418 17276 14424
rect 17052 13462 17080 14418
rect 17868 14408 17920 14414
rect 17868 14350 17920 14356
rect 17132 14068 17184 14074
rect 17132 14010 17184 14016
rect 17040 13456 17092 13462
rect 17040 13398 17092 13404
rect 17040 12640 17092 12646
rect 17040 12582 17092 12588
rect 16948 12164 17000 12170
rect 16948 12106 17000 12112
rect 17052 12073 17080 12582
rect 17038 12064 17094 12073
rect 17038 11999 17094 12008
rect 17052 11626 17080 11999
rect 17040 11620 17092 11626
rect 17040 11562 17092 11568
rect 16948 11552 17000 11558
rect 16948 11494 17000 11500
rect 16960 11218 16988 11494
rect 16948 11212 17000 11218
rect 16948 11154 17000 11160
rect 17144 10146 17172 14010
rect 17776 13864 17828 13870
rect 17776 13806 17828 13812
rect 17788 12986 17816 13806
rect 17880 13682 17908 14350
rect 17972 13870 18000 15982
rect 18156 15910 18184 19654
rect 18236 16176 18288 16182
rect 18236 16118 18288 16124
rect 18144 15904 18196 15910
rect 18144 15846 18196 15852
rect 18144 15020 18196 15026
rect 18144 14962 18196 14968
rect 18050 13968 18106 13977
rect 18050 13903 18106 13912
rect 17960 13864 18012 13870
rect 17960 13806 18012 13812
rect 18064 13734 18092 13903
rect 18052 13728 18104 13734
rect 17880 13654 18000 13682
rect 18052 13670 18104 13676
rect 17972 13394 18000 13654
rect 17960 13388 18012 13394
rect 17960 13330 18012 13336
rect 17776 12980 17828 12986
rect 17776 12922 17828 12928
rect 17684 12368 17736 12374
rect 17684 12310 17736 12316
rect 17224 11756 17276 11762
rect 17224 11698 17276 11704
rect 17236 11354 17264 11698
rect 17224 11348 17276 11354
rect 17224 11290 17276 11296
rect 17236 10674 17264 11290
rect 17696 11286 17724 12310
rect 17684 11280 17736 11286
rect 17684 11222 17736 11228
rect 17592 11008 17644 11014
rect 17592 10950 17644 10956
rect 17498 10704 17554 10713
rect 17224 10668 17276 10674
rect 17604 10674 17632 10950
rect 17498 10639 17500 10648
rect 17224 10610 17276 10616
rect 17552 10639 17554 10648
rect 17592 10668 17644 10674
rect 17500 10610 17552 10616
rect 17592 10610 17644 10616
rect 17776 10668 17828 10674
rect 17776 10610 17828 10616
rect 17868 10668 17920 10674
rect 17920 10628 18000 10656
rect 17868 10610 17920 10616
rect 17052 10118 17172 10146
rect 17236 10130 17264 10610
rect 17788 10198 17816 10610
rect 17776 10192 17828 10198
rect 17776 10134 17828 10140
rect 17224 10124 17276 10130
rect 16948 10056 17000 10062
rect 16946 10024 16948 10033
rect 17000 10024 17002 10033
rect 16946 9959 17002 9968
rect 16856 8492 16908 8498
rect 16856 8434 16908 8440
rect 16764 8288 16816 8294
rect 16764 8230 16816 8236
rect 16580 7812 16632 7818
rect 16580 7754 16632 7760
rect 16592 7585 16620 7754
rect 16672 7744 16724 7750
rect 16672 7686 16724 7692
rect 16578 7576 16634 7585
rect 16578 7511 16634 7520
rect 16580 7404 16632 7410
rect 16580 7346 16632 7352
rect 16592 7313 16620 7346
rect 16578 7304 16634 7313
rect 16578 7239 16634 7248
rect 16684 7002 16712 7686
rect 16776 7410 16804 8230
rect 16948 8016 17000 8022
rect 16868 7976 16948 8004
rect 16764 7404 16816 7410
rect 16764 7346 16816 7352
rect 16868 7274 16896 7976
rect 16948 7958 17000 7964
rect 17052 7886 17080 10118
rect 17224 10066 17276 10072
rect 17408 10124 17460 10130
rect 17408 10066 17460 10072
rect 17420 9994 17448 10066
rect 17972 10033 18000 10628
rect 17958 10024 18014 10033
rect 17408 9988 17460 9994
rect 17958 9959 18014 9968
rect 17408 9930 17460 9936
rect 17316 9104 17368 9110
rect 17316 9046 17368 9052
rect 17132 8832 17184 8838
rect 17132 8774 17184 8780
rect 17144 8498 17172 8774
rect 17328 8566 17356 9046
rect 17316 8560 17368 8566
rect 17316 8502 17368 8508
rect 17132 8492 17184 8498
rect 17132 8434 17184 8440
rect 17222 8256 17278 8265
rect 17222 8191 17278 8200
rect 17236 8090 17264 8191
rect 17224 8084 17276 8090
rect 17224 8026 17276 8032
rect 17130 7984 17186 7993
rect 17420 7970 17448 9930
rect 17868 9376 17920 9382
rect 17868 9318 17920 9324
rect 17592 8832 17644 8838
rect 17592 8774 17644 8780
rect 17130 7919 17186 7928
rect 17236 7942 17448 7970
rect 17144 7886 17172 7919
rect 16948 7880 17000 7886
rect 16948 7822 17000 7828
rect 17040 7880 17092 7886
rect 17040 7822 17092 7828
rect 17132 7880 17184 7886
rect 17132 7822 17184 7828
rect 16960 7290 16988 7822
rect 17040 7744 17092 7750
rect 17040 7686 17092 7692
rect 17052 7410 17080 7686
rect 17236 7426 17264 7942
rect 17604 7886 17632 8774
rect 17684 7948 17736 7954
rect 17684 7890 17736 7896
rect 17592 7880 17644 7886
rect 17512 7840 17592 7868
rect 17408 7744 17460 7750
rect 17408 7686 17460 7692
rect 17040 7404 17092 7410
rect 17236 7398 17356 7426
rect 17420 7410 17448 7686
rect 17040 7346 17092 7352
rect 17328 7342 17356 7398
rect 17408 7404 17460 7410
rect 17408 7346 17460 7352
rect 17316 7336 17368 7342
rect 16960 7274 17080 7290
rect 17316 7278 17368 7284
rect 16856 7268 16908 7274
rect 16960 7268 17092 7274
rect 16960 7262 17040 7268
rect 16856 7210 16908 7216
rect 17040 7210 17092 7216
rect 16672 6996 16724 7002
rect 16672 6938 16724 6944
rect 16488 6792 16540 6798
rect 16488 6734 16540 6740
rect 16304 6656 16356 6662
rect 16304 6598 16356 6604
rect 16028 6384 16080 6390
rect 16028 6326 16080 6332
rect 16500 6322 16528 6734
rect 17052 6390 17080 7210
rect 17328 7002 17356 7278
rect 17512 7177 17540 7840
rect 17592 7822 17644 7828
rect 17696 7546 17724 7890
rect 17776 7880 17828 7886
rect 17774 7848 17776 7857
rect 17828 7848 17830 7857
rect 17774 7783 17830 7792
rect 17684 7540 17736 7546
rect 17684 7482 17736 7488
rect 17880 7410 17908 9318
rect 17972 8906 18000 9959
rect 17960 8900 18012 8906
rect 17960 8842 18012 8848
rect 17972 7410 18000 8842
rect 18064 7970 18092 13670
rect 18156 10810 18184 14962
rect 18248 14346 18276 16118
rect 18340 16046 18368 20810
rect 18696 20800 18748 20806
rect 18696 20742 18748 20748
rect 18512 20528 18564 20534
rect 18564 20488 18644 20516
rect 18512 20470 18564 20476
rect 18512 20256 18564 20262
rect 18512 20198 18564 20204
rect 18524 19514 18552 20198
rect 18512 19508 18564 19514
rect 18512 19450 18564 19456
rect 18616 19334 18644 20488
rect 18708 19378 18736 20742
rect 18800 19854 18828 22066
rect 18788 19848 18840 19854
rect 18788 19790 18840 19796
rect 18800 19514 18828 19790
rect 18892 19786 18920 23666
rect 19076 22094 19104 24210
rect 18984 22066 19104 22094
rect 18984 19922 19012 22066
rect 19064 21548 19116 21554
rect 19064 21490 19116 21496
rect 19076 21146 19104 21490
rect 19064 21140 19116 21146
rect 19064 21082 19116 21088
rect 19064 20936 19116 20942
rect 19064 20878 19116 20884
rect 18972 19916 19024 19922
rect 18972 19858 19024 19864
rect 18880 19780 18932 19786
rect 18880 19722 18932 19728
rect 18788 19508 18840 19514
rect 18788 19450 18840 19456
rect 18524 19306 18644 19334
rect 18696 19372 18748 19378
rect 18696 19314 18748 19320
rect 18524 18766 18552 19306
rect 18892 19174 18920 19722
rect 18880 19168 18932 19174
rect 18880 19110 18932 19116
rect 18512 18760 18564 18766
rect 18512 18702 18564 18708
rect 18420 17672 18472 17678
rect 18420 17614 18472 17620
rect 18328 16040 18380 16046
rect 18328 15982 18380 15988
rect 18328 14952 18380 14958
rect 18328 14894 18380 14900
rect 18236 14340 18288 14346
rect 18236 14282 18288 14288
rect 18236 14000 18288 14006
rect 18236 13942 18288 13948
rect 18144 10804 18196 10810
rect 18144 10746 18196 10752
rect 18144 10668 18196 10674
rect 18144 10610 18196 10616
rect 18156 10130 18184 10610
rect 18144 10124 18196 10130
rect 18144 10066 18196 10072
rect 18144 9580 18196 9586
rect 18144 9522 18196 9528
rect 18156 8430 18184 9522
rect 18248 9518 18276 13942
rect 18340 11150 18368 14894
rect 18432 14414 18460 17614
rect 18524 16250 18552 18702
rect 18788 18420 18840 18426
rect 18788 18362 18840 18368
rect 18800 17678 18828 18362
rect 18788 17672 18840 17678
rect 18788 17614 18840 17620
rect 18604 17536 18656 17542
rect 18604 17478 18656 17484
rect 18788 17536 18840 17542
rect 18788 17478 18840 17484
rect 18616 17338 18644 17478
rect 18604 17332 18656 17338
rect 18604 17274 18656 17280
rect 18616 16726 18644 17274
rect 18800 16794 18828 17478
rect 18788 16788 18840 16794
rect 18788 16730 18840 16736
rect 18604 16720 18656 16726
rect 18604 16662 18656 16668
rect 18696 16584 18748 16590
rect 18696 16526 18748 16532
rect 18512 16244 18564 16250
rect 18512 16186 18564 16192
rect 18708 16182 18736 16526
rect 18788 16244 18840 16250
rect 18788 16186 18840 16192
rect 18696 16176 18748 16182
rect 18696 16118 18748 16124
rect 18512 16108 18564 16114
rect 18512 16050 18564 16056
rect 18524 15162 18552 16050
rect 18696 15972 18748 15978
rect 18696 15914 18748 15920
rect 18604 15904 18656 15910
rect 18604 15846 18656 15852
rect 18616 15366 18644 15846
rect 18708 15706 18736 15914
rect 18696 15700 18748 15706
rect 18696 15642 18748 15648
rect 18604 15360 18656 15366
rect 18604 15302 18656 15308
rect 18512 15156 18564 15162
rect 18512 15098 18564 15104
rect 18616 15042 18644 15302
rect 18524 15014 18644 15042
rect 18420 14408 18472 14414
rect 18420 14350 18472 14356
rect 18420 14000 18472 14006
rect 18420 13942 18472 13948
rect 18432 13326 18460 13942
rect 18420 13320 18472 13326
rect 18420 13262 18472 13268
rect 18524 12850 18552 15014
rect 18800 14090 18828 16186
rect 18604 14068 18656 14074
rect 18604 14010 18656 14016
rect 18708 14062 18828 14090
rect 18616 13802 18644 14010
rect 18604 13796 18656 13802
rect 18604 13738 18656 13744
rect 18708 13258 18736 14062
rect 18892 14006 18920 19110
rect 18880 14000 18932 14006
rect 18880 13942 18932 13948
rect 18984 13938 19012 19858
rect 19076 19446 19104 20878
rect 19156 20868 19208 20874
rect 19156 20810 19208 20816
rect 19168 20466 19196 20810
rect 19260 20788 19288 24210
rect 20640 24206 20668 24754
rect 21744 24410 21772 24754
rect 21836 24410 21864 25230
rect 22192 25220 22244 25226
rect 22192 25162 22244 25168
rect 22204 24750 22232 25162
rect 22192 24744 22244 24750
rect 22192 24686 22244 24692
rect 21916 24676 21968 24682
rect 21916 24618 21968 24624
rect 22008 24676 22060 24682
rect 22008 24618 22060 24624
rect 21732 24404 21784 24410
rect 21732 24346 21784 24352
rect 21824 24404 21876 24410
rect 21824 24346 21876 24352
rect 21928 24274 21956 24618
rect 22020 24410 22048 24618
rect 22008 24404 22060 24410
rect 22008 24346 22060 24352
rect 21916 24268 21968 24274
rect 21744 24228 21916 24256
rect 20628 24200 20680 24206
rect 20628 24142 20680 24148
rect 21548 24200 21600 24206
rect 21548 24142 21600 24148
rect 19432 23724 19484 23730
rect 19432 23666 19484 23672
rect 19616 23724 19668 23730
rect 19616 23666 19668 23672
rect 20444 23724 20496 23730
rect 20444 23666 20496 23672
rect 19444 23254 19472 23666
rect 19628 23322 19656 23666
rect 19616 23316 19668 23322
rect 19616 23258 19668 23264
rect 19340 23248 19392 23254
rect 19340 23190 19392 23196
rect 19432 23248 19484 23254
rect 19432 23190 19484 23196
rect 19352 23050 19380 23190
rect 20456 23118 20484 23666
rect 20352 23112 20404 23118
rect 20352 23054 20404 23060
rect 20444 23112 20496 23118
rect 20444 23054 20496 23060
rect 19340 23044 19392 23050
rect 19340 22986 19392 22992
rect 19432 22976 19484 22982
rect 19432 22918 19484 22924
rect 19444 22778 19472 22918
rect 19432 22772 19484 22778
rect 19432 22714 19484 22720
rect 19616 22432 19668 22438
rect 19616 22374 19668 22380
rect 19432 21480 19484 21486
rect 19432 21422 19484 21428
rect 19260 20760 19380 20788
rect 19156 20460 19208 20466
rect 19156 20402 19208 20408
rect 19248 20392 19300 20398
rect 19154 20360 19210 20369
rect 19352 20380 19380 20760
rect 19300 20352 19380 20380
rect 19248 20334 19300 20340
rect 19154 20295 19156 20304
rect 19208 20295 19210 20304
rect 19156 20266 19208 20272
rect 19064 19440 19116 19446
rect 19064 19382 19116 19388
rect 19260 18970 19288 20334
rect 19340 19984 19392 19990
rect 19340 19926 19392 19932
rect 19352 19446 19380 19926
rect 19340 19440 19392 19446
rect 19340 19382 19392 19388
rect 19248 18964 19300 18970
rect 19248 18906 19300 18912
rect 19340 18692 19392 18698
rect 19340 18634 19392 18640
rect 19248 17672 19300 17678
rect 19062 17640 19118 17649
rect 19248 17614 19300 17620
rect 19062 17575 19118 17584
rect 19156 17604 19208 17610
rect 19076 17202 19104 17575
rect 19156 17546 19208 17552
rect 19064 17196 19116 17202
rect 19064 17138 19116 17144
rect 19076 17105 19104 17138
rect 19062 17096 19118 17105
rect 19062 17031 19118 17040
rect 19064 16584 19116 16590
rect 19064 16526 19116 16532
rect 19076 16250 19104 16526
rect 19064 16244 19116 16250
rect 19064 16186 19116 16192
rect 19168 14482 19196 17546
rect 19260 16658 19288 17614
rect 19248 16652 19300 16658
rect 19248 16594 19300 16600
rect 19352 15910 19380 18634
rect 19340 15904 19392 15910
rect 19340 15846 19392 15852
rect 19156 14476 19208 14482
rect 19156 14418 19208 14424
rect 19064 14408 19116 14414
rect 19064 14350 19116 14356
rect 18788 13932 18840 13938
rect 18788 13874 18840 13880
rect 18972 13932 19024 13938
rect 18972 13874 19024 13880
rect 18696 13252 18748 13258
rect 18696 13194 18748 13200
rect 18696 12980 18748 12986
rect 18800 12968 18828 13874
rect 18880 13864 18932 13870
rect 18880 13806 18932 13812
rect 18892 13394 18920 13806
rect 18972 13728 19024 13734
rect 18972 13670 19024 13676
rect 18984 13530 19012 13670
rect 18972 13524 19024 13530
rect 18972 13466 19024 13472
rect 18880 13388 18932 13394
rect 18880 13330 18932 13336
rect 18748 12940 18828 12968
rect 18696 12922 18748 12928
rect 18512 12844 18564 12850
rect 18512 12786 18564 12792
rect 18708 12374 18736 12922
rect 19076 12434 19104 14350
rect 19168 14006 19196 14418
rect 19156 14000 19208 14006
rect 19156 13942 19208 13948
rect 19076 12406 19196 12434
rect 18696 12368 18748 12374
rect 18696 12310 18748 12316
rect 18420 12096 18472 12102
rect 18420 12038 18472 12044
rect 18432 11762 18460 12038
rect 18420 11756 18472 11762
rect 18420 11698 18472 11704
rect 18604 11552 18656 11558
rect 18604 11494 18656 11500
rect 18788 11552 18840 11558
rect 18788 11494 18840 11500
rect 18328 11144 18380 11150
rect 18328 11086 18380 11092
rect 18340 10198 18368 11086
rect 18512 11076 18564 11082
rect 18512 11018 18564 11024
rect 18420 10804 18472 10810
rect 18420 10746 18472 10752
rect 18328 10192 18380 10198
rect 18328 10134 18380 10140
rect 18328 10056 18380 10062
rect 18326 10024 18328 10033
rect 18380 10024 18382 10033
rect 18326 9959 18382 9968
rect 18236 9512 18288 9518
rect 18236 9454 18288 9460
rect 18248 9178 18276 9454
rect 18236 9172 18288 9178
rect 18236 9114 18288 9120
rect 18432 8838 18460 10746
rect 18524 10742 18552 11018
rect 18512 10736 18564 10742
rect 18512 10678 18564 10684
rect 18616 10538 18644 11494
rect 18696 11348 18748 11354
rect 18696 11290 18748 11296
rect 18604 10532 18656 10538
rect 18604 10474 18656 10480
rect 18420 8832 18472 8838
rect 18420 8774 18472 8780
rect 18144 8424 18196 8430
rect 18144 8366 18196 8372
rect 18512 8424 18564 8430
rect 18512 8366 18564 8372
rect 18064 7942 18184 7970
rect 18052 7812 18104 7818
rect 18052 7754 18104 7760
rect 18064 7546 18092 7754
rect 18156 7546 18184 7942
rect 18524 7886 18552 8366
rect 18616 7886 18644 10474
rect 18420 7880 18472 7886
rect 18420 7822 18472 7828
rect 18512 7880 18564 7886
rect 18604 7880 18656 7886
rect 18512 7822 18564 7828
rect 18602 7848 18604 7857
rect 18656 7848 18658 7857
rect 18236 7812 18288 7818
rect 18236 7754 18288 7760
rect 18052 7540 18104 7546
rect 18052 7482 18104 7488
rect 18144 7540 18196 7546
rect 18144 7482 18196 7488
rect 17592 7404 17644 7410
rect 17592 7346 17644 7352
rect 17868 7404 17920 7410
rect 17868 7346 17920 7352
rect 17960 7404 18012 7410
rect 17960 7346 18012 7352
rect 17498 7168 17554 7177
rect 17498 7103 17554 7112
rect 17604 7002 17632 7346
rect 17316 6996 17368 7002
rect 17316 6938 17368 6944
rect 17592 6996 17644 7002
rect 17592 6938 17644 6944
rect 18156 6866 18184 7482
rect 18248 7410 18276 7754
rect 18432 7546 18460 7822
rect 18420 7540 18472 7546
rect 18420 7482 18472 7488
rect 18524 7478 18552 7822
rect 18602 7783 18658 7792
rect 18512 7472 18564 7478
rect 18512 7414 18564 7420
rect 18236 7404 18288 7410
rect 18236 7346 18288 7352
rect 18604 7336 18656 7342
rect 18604 7278 18656 7284
rect 18144 6860 18196 6866
rect 18144 6802 18196 6808
rect 18616 6458 18644 7278
rect 18708 6798 18736 11290
rect 18800 10810 18828 11494
rect 18972 11076 19024 11082
rect 18972 11018 19024 11024
rect 18788 10804 18840 10810
rect 18788 10746 18840 10752
rect 18788 10056 18840 10062
rect 18788 9998 18840 10004
rect 18800 9722 18828 9998
rect 18788 9716 18840 9722
rect 18788 9658 18840 9664
rect 18880 9512 18932 9518
rect 18880 9454 18932 9460
rect 18892 9330 18920 9454
rect 18984 9450 19012 11018
rect 19064 9988 19116 9994
rect 19064 9930 19116 9936
rect 19076 9654 19104 9930
rect 19064 9648 19116 9654
rect 19064 9590 19116 9596
rect 18972 9444 19024 9450
rect 18972 9386 19024 9392
rect 18892 9302 19012 9330
rect 18788 8832 18840 8838
rect 18788 8774 18840 8780
rect 18800 7886 18828 8774
rect 18984 8498 19012 9302
rect 18972 8492 19024 8498
rect 18972 8434 19024 8440
rect 18878 7984 18934 7993
rect 18878 7919 18934 7928
rect 18892 7886 18920 7919
rect 18788 7880 18840 7886
rect 18788 7822 18840 7828
rect 18880 7880 18932 7886
rect 18880 7822 18932 7828
rect 18800 7449 18828 7822
rect 18786 7440 18842 7449
rect 18786 7375 18842 7384
rect 18984 6866 19012 8434
rect 19168 7818 19196 12406
rect 19352 12238 19380 15846
rect 19444 15638 19472 21422
rect 19524 21344 19576 21350
rect 19524 21286 19576 21292
rect 19536 21078 19564 21286
rect 19628 21078 19656 22374
rect 19708 21684 19760 21690
rect 19708 21626 19760 21632
rect 19524 21072 19576 21078
rect 19524 21014 19576 21020
rect 19616 21072 19668 21078
rect 19616 21014 19668 21020
rect 19616 20936 19668 20942
rect 19720 20924 19748 21626
rect 20364 21622 20392 23054
rect 20456 22710 20484 23054
rect 20444 22704 20496 22710
rect 20444 22646 20496 22652
rect 20536 22568 20588 22574
rect 20536 22510 20588 22516
rect 19984 21616 20036 21622
rect 19984 21558 20036 21564
rect 20352 21616 20404 21622
rect 20352 21558 20404 21564
rect 19800 21344 19852 21350
rect 19798 21312 19800 21321
rect 19852 21312 19854 21321
rect 19798 21247 19854 21256
rect 19668 20896 19748 20924
rect 19616 20878 19668 20884
rect 19524 20800 19576 20806
rect 19524 20742 19576 20748
rect 19536 20534 19564 20742
rect 19616 20596 19668 20602
rect 19616 20538 19668 20544
rect 19892 20596 19944 20602
rect 19996 20584 20024 21558
rect 20548 20942 20576 22510
rect 20076 20936 20128 20942
rect 20076 20878 20128 20884
rect 20168 20936 20220 20942
rect 20168 20878 20220 20884
rect 20536 20936 20588 20942
rect 20536 20878 20588 20884
rect 19944 20556 20024 20584
rect 19892 20538 19944 20544
rect 19524 20528 19576 20534
rect 19524 20470 19576 20476
rect 19524 19780 19576 19786
rect 19628 19768 19656 20538
rect 19892 20256 19944 20262
rect 19892 20198 19944 20204
rect 19904 19922 19932 20198
rect 19892 19916 19944 19922
rect 19892 19858 19944 19864
rect 19996 19854 20024 20556
rect 20088 20262 20116 20878
rect 20076 20256 20128 20262
rect 20076 20198 20128 20204
rect 19708 19848 19760 19854
rect 19708 19790 19760 19796
rect 19984 19848 20036 19854
rect 19984 19790 20036 19796
rect 19576 19740 19656 19768
rect 19524 19722 19576 19728
rect 19536 19242 19564 19722
rect 19720 19446 19748 19790
rect 20088 19718 20116 20198
rect 20180 19990 20208 20878
rect 20260 20868 20312 20874
rect 20260 20810 20312 20816
rect 20168 19984 20220 19990
rect 20168 19926 20220 19932
rect 20272 19854 20300 20810
rect 20352 20800 20404 20806
rect 20352 20742 20404 20748
rect 20364 19922 20392 20742
rect 20640 20466 20668 24142
rect 21560 23866 21588 24142
rect 21548 23860 21600 23866
rect 21548 23802 21600 23808
rect 21744 23730 21772 24228
rect 21916 24210 21968 24216
rect 22480 24256 22508 26250
rect 23032 25498 23060 26250
rect 23768 25770 23796 27338
rect 24228 27130 24256 27406
rect 24216 27124 24268 27130
rect 24216 27066 24268 27072
rect 24412 26994 24440 27406
rect 24596 27033 24624 27526
rect 24860 27474 24912 27480
rect 24676 27464 24728 27470
rect 24676 27406 24728 27412
rect 24582 27024 24638 27033
rect 24400 26988 24452 26994
rect 24688 26994 24716 27406
rect 24768 27124 24820 27130
rect 24768 27066 24820 27072
rect 24780 26994 24808 27066
rect 24582 26959 24638 26968
rect 24676 26988 24728 26994
rect 24400 26930 24452 26936
rect 24492 26920 24544 26926
rect 24492 26862 24544 26868
rect 24216 26784 24268 26790
rect 24216 26726 24268 26732
rect 24228 26586 24256 26726
rect 24216 26580 24268 26586
rect 24216 26522 24268 26528
rect 24228 26382 24256 26522
rect 24216 26376 24268 26382
rect 24216 26318 24268 26324
rect 23756 25764 23808 25770
rect 23756 25706 23808 25712
rect 23020 25492 23072 25498
rect 23020 25434 23072 25440
rect 22744 25424 22796 25430
rect 22744 25366 22796 25372
rect 22652 25288 22704 25294
rect 22652 25230 22704 25236
rect 22664 24886 22692 25230
rect 22652 24880 22704 24886
rect 22652 24822 22704 24828
rect 22560 24268 22612 24274
rect 22480 24228 22560 24256
rect 22192 24132 22244 24138
rect 22192 24074 22244 24080
rect 21824 24064 21876 24070
rect 21824 24006 21876 24012
rect 21836 23746 21864 24006
rect 22008 23792 22060 23798
rect 21836 23740 22008 23746
rect 21836 23734 22060 23740
rect 21732 23724 21784 23730
rect 21836 23718 22048 23734
rect 21732 23666 21784 23672
rect 22204 23322 22232 24074
rect 22192 23316 22244 23322
rect 22192 23258 22244 23264
rect 20812 23112 20864 23118
rect 20812 23054 20864 23060
rect 20824 22778 20852 23054
rect 22480 23050 22508 24228
rect 22560 24210 22612 24216
rect 22756 23118 22784 25366
rect 23296 25356 23348 25362
rect 23296 25298 23348 25304
rect 23020 25220 23072 25226
rect 23020 25162 23072 25168
rect 23032 25106 23060 25162
rect 23032 25078 23152 25106
rect 23124 23662 23152 25078
rect 23308 24410 23336 25298
rect 23388 25288 23440 25294
rect 23388 25230 23440 25236
rect 23296 24404 23348 24410
rect 23296 24346 23348 24352
rect 23400 23730 23428 25230
rect 23572 25220 23624 25226
rect 23572 25162 23624 25168
rect 23480 24132 23532 24138
rect 23480 24074 23532 24080
rect 23492 23798 23520 24074
rect 23480 23792 23532 23798
rect 23480 23734 23532 23740
rect 23388 23724 23440 23730
rect 23388 23666 23440 23672
rect 23112 23656 23164 23662
rect 23112 23598 23164 23604
rect 23400 23322 23428 23666
rect 23584 23594 23612 25162
rect 23664 25152 23716 25158
rect 23664 25094 23716 25100
rect 23676 24070 23704 25094
rect 23848 24744 23900 24750
rect 23848 24686 23900 24692
rect 23664 24064 23716 24070
rect 23664 24006 23716 24012
rect 23572 23588 23624 23594
rect 23572 23530 23624 23536
rect 23480 23520 23532 23526
rect 23480 23462 23532 23468
rect 23388 23316 23440 23322
rect 23388 23258 23440 23264
rect 23492 23186 23520 23462
rect 23676 23254 23704 24006
rect 23664 23248 23716 23254
rect 23664 23190 23716 23196
rect 23480 23180 23532 23186
rect 23480 23122 23532 23128
rect 23860 23118 23888 24686
rect 24308 24200 24360 24206
rect 24136 24148 24308 24154
rect 24136 24142 24360 24148
rect 24136 24138 24348 24142
rect 24124 24132 24348 24138
rect 24176 24126 24348 24132
rect 24124 24074 24176 24080
rect 24504 24052 24532 26862
rect 24596 26246 24624 26959
rect 24676 26930 24728 26936
rect 24768 26988 24820 26994
rect 24768 26930 24820 26936
rect 24688 26314 24716 26930
rect 24872 26586 24900 27474
rect 24964 27033 24992 28018
rect 25056 27674 25084 28018
rect 25412 28008 25464 28014
rect 25412 27950 25464 27956
rect 25044 27668 25096 27674
rect 25044 27610 25096 27616
rect 24950 27024 25006 27033
rect 24950 26959 24952 26968
rect 25004 26959 25006 26968
rect 25056 26976 25084 27610
rect 25318 27568 25374 27577
rect 25240 27512 25318 27520
rect 25240 27492 25320 27512
rect 25136 26988 25188 26994
rect 25056 26948 25136 26976
rect 24952 26930 25004 26936
rect 25136 26930 25188 26936
rect 25240 26926 25268 27492
rect 25372 27503 25374 27512
rect 25320 27474 25372 27480
rect 25424 27062 25452 27950
rect 25780 27600 25832 27606
rect 25780 27542 25832 27548
rect 25792 27470 25820 27542
rect 25504 27464 25556 27470
rect 25504 27406 25556 27412
rect 25780 27464 25832 27470
rect 25780 27406 25832 27412
rect 25412 27056 25464 27062
rect 25412 26998 25464 27004
rect 25228 26920 25280 26926
rect 25228 26862 25280 26868
rect 24860 26580 24912 26586
rect 24860 26522 24912 26528
rect 24952 26512 25004 26518
rect 24952 26454 25004 26460
rect 24860 26376 24912 26382
rect 24860 26318 24912 26324
rect 24676 26308 24728 26314
rect 24676 26250 24728 26256
rect 24584 26240 24636 26246
rect 24584 26182 24636 26188
rect 24768 25220 24820 25226
rect 24768 25162 24820 25168
rect 24780 24818 24808 25162
rect 24768 24812 24820 24818
rect 24768 24754 24820 24760
rect 24676 24200 24728 24206
rect 24676 24142 24728 24148
rect 24584 24064 24636 24070
rect 24504 24024 24584 24052
rect 24584 24006 24636 24012
rect 24032 23724 24084 23730
rect 24032 23666 24084 23672
rect 24044 23118 24072 23666
rect 24216 23520 24268 23526
rect 24216 23462 24268 23468
rect 24228 23118 24256 23462
rect 24400 23180 24452 23186
rect 24400 23122 24452 23128
rect 22744 23112 22796 23118
rect 22744 23054 22796 23060
rect 23848 23112 23900 23118
rect 23848 23054 23900 23060
rect 24032 23112 24084 23118
rect 24032 23054 24084 23060
rect 24216 23112 24268 23118
rect 24216 23054 24268 23060
rect 22468 23044 22520 23050
rect 22468 22986 22520 22992
rect 20812 22772 20864 22778
rect 20812 22714 20864 22720
rect 20996 22636 21048 22642
rect 20996 22578 21048 22584
rect 22284 22636 22336 22642
rect 22284 22578 22336 22584
rect 21008 22234 21036 22578
rect 20996 22228 21048 22234
rect 20996 22170 21048 22176
rect 21548 22228 21600 22234
rect 21548 22170 21600 22176
rect 21088 21548 21140 21554
rect 21088 21490 21140 21496
rect 21100 20942 21128 21490
rect 21180 21412 21232 21418
rect 21180 21354 21232 21360
rect 21192 21146 21220 21354
rect 21364 21344 21416 21350
rect 21364 21286 21416 21292
rect 21180 21140 21232 21146
rect 21180 21082 21232 21088
rect 21088 20936 21140 20942
rect 21088 20878 21140 20884
rect 20904 20800 20956 20806
rect 20904 20742 20956 20748
rect 20628 20460 20680 20466
rect 20628 20402 20680 20408
rect 20640 20330 20668 20402
rect 20628 20324 20680 20330
rect 20628 20266 20680 20272
rect 20352 19916 20404 19922
rect 20352 19858 20404 19864
rect 20260 19848 20312 19854
rect 20260 19790 20312 19796
rect 20076 19712 20128 19718
rect 20076 19654 20128 19660
rect 19708 19440 19760 19446
rect 19708 19382 19760 19388
rect 19720 19334 19748 19382
rect 20088 19378 20116 19654
rect 19628 19306 19748 19334
rect 20076 19372 20128 19378
rect 20076 19314 20128 19320
rect 19524 19236 19576 19242
rect 19524 19178 19576 19184
rect 19536 16726 19564 19178
rect 19628 17626 19656 19306
rect 19708 19168 19760 19174
rect 19708 19110 19760 19116
rect 19720 17746 19748 19110
rect 19800 17808 19852 17814
rect 19800 17750 19852 17756
rect 20628 17808 20680 17814
rect 20628 17750 20680 17756
rect 19708 17740 19760 17746
rect 19708 17682 19760 17688
rect 19628 17598 19748 17626
rect 19524 16720 19576 16726
rect 19524 16662 19576 16668
rect 19432 15632 19484 15638
rect 19432 15574 19484 15580
rect 19432 15496 19484 15502
rect 19432 15438 19484 15444
rect 19444 12442 19472 15438
rect 19536 13841 19564 16662
rect 19720 16454 19748 17598
rect 19812 16794 19840 17750
rect 20260 17536 20312 17542
rect 20260 17478 20312 17484
rect 20272 17202 20300 17478
rect 20534 17368 20590 17377
rect 20534 17303 20536 17312
rect 20588 17303 20590 17312
rect 20536 17274 20588 17280
rect 20640 17202 20668 17750
rect 20916 17746 20944 20742
rect 21100 20602 21128 20878
rect 21088 20596 21140 20602
rect 21088 20538 21140 20544
rect 21192 20466 21220 21082
rect 21376 21078 21404 21286
rect 21364 21072 21416 21078
rect 21364 21014 21416 21020
rect 21376 20466 21404 21014
rect 21560 21010 21588 22170
rect 22192 21480 22244 21486
rect 22192 21422 22244 21428
rect 22008 21072 22060 21078
rect 22008 21014 22060 21020
rect 21548 21004 21600 21010
rect 21548 20946 21600 20952
rect 21180 20460 21232 20466
rect 21180 20402 21232 20408
rect 21364 20460 21416 20466
rect 21364 20402 21416 20408
rect 21560 19854 21588 20946
rect 21916 20800 21968 20806
rect 21916 20742 21968 20748
rect 21824 20528 21876 20534
rect 21824 20470 21876 20476
rect 21548 19848 21600 19854
rect 21548 19790 21600 19796
rect 21836 19786 21864 20470
rect 21928 20262 21956 20742
rect 22020 20602 22048 21014
rect 22204 20942 22232 21422
rect 22100 20936 22152 20942
rect 22100 20878 22152 20884
rect 22192 20936 22244 20942
rect 22192 20878 22244 20884
rect 22008 20596 22060 20602
rect 22008 20538 22060 20544
rect 21916 20256 21968 20262
rect 21916 20198 21968 20204
rect 21928 19854 21956 20198
rect 22020 19854 22048 20538
rect 22112 19990 22140 20878
rect 22296 20874 22324 22578
rect 23296 21684 23348 21690
rect 23296 21626 23348 21632
rect 23112 21548 23164 21554
rect 23112 21490 23164 21496
rect 22928 21480 22980 21486
rect 22928 21422 22980 21428
rect 22744 21412 22796 21418
rect 22744 21354 22796 21360
rect 22560 21004 22612 21010
rect 22480 20964 22560 20992
rect 22376 20936 22428 20942
rect 22376 20878 22428 20884
rect 22284 20868 22336 20874
rect 22284 20810 22336 20816
rect 22388 20806 22416 20878
rect 22192 20800 22244 20806
rect 22192 20742 22244 20748
rect 22376 20800 22428 20806
rect 22376 20742 22428 20748
rect 22204 20602 22232 20742
rect 22192 20596 22244 20602
rect 22192 20538 22244 20544
rect 22100 19984 22152 19990
rect 22100 19926 22152 19932
rect 22204 19854 22232 20538
rect 22480 19854 22508 20964
rect 22560 20946 22612 20952
rect 22756 20942 22784 21354
rect 22744 20936 22796 20942
rect 22744 20878 22796 20884
rect 22744 20800 22796 20806
rect 22744 20742 22796 20748
rect 22560 20392 22612 20398
rect 22756 20369 22784 20742
rect 22836 20528 22888 20534
rect 22836 20470 22888 20476
rect 22560 20334 22612 20340
rect 22742 20360 22798 20369
rect 22572 20058 22600 20334
rect 22742 20295 22798 20304
rect 22560 20052 22612 20058
rect 22560 19994 22612 20000
rect 22652 19916 22704 19922
rect 22652 19858 22704 19864
rect 21916 19848 21968 19854
rect 21916 19790 21968 19796
rect 22008 19848 22060 19854
rect 22008 19790 22060 19796
rect 22192 19848 22244 19854
rect 22192 19790 22244 19796
rect 22468 19848 22520 19854
rect 22468 19790 22520 19796
rect 22560 19848 22612 19854
rect 22560 19790 22612 19796
rect 21824 19780 21876 19786
rect 21824 19722 21876 19728
rect 22376 19780 22428 19786
rect 22376 19722 22428 19728
rect 22100 19712 22152 19718
rect 22100 19654 22152 19660
rect 22192 19712 22244 19718
rect 22244 19672 22324 19700
rect 22192 19654 22244 19660
rect 22112 19514 22140 19654
rect 22100 19508 22152 19514
rect 22100 19450 22152 19456
rect 21916 18216 21968 18222
rect 21916 18158 21968 18164
rect 20904 17740 20956 17746
rect 20904 17682 20956 17688
rect 20812 17672 20864 17678
rect 20812 17614 20864 17620
rect 20720 17536 20772 17542
rect 20720 17478 20772 17484
rect 20260 17196 20312 17202
rect 20260 17138 20312 17144
rect 20352 17196 20404 17202
rect 20352 17138 20404 17144
rect 20628 17196 20680 17202
rect 20628 17138 20680 17144
rect 19892 16992 19944 16998
rect 19892 16934 19944 16940
rect 19800 16788 19852 16794
rect 19800 16730 19852 16736
rect 19708 16448 19760 16454
rect 19708 16390 19760 16396
rect 19616 15564 19668 15570
rect 19616 15506 19668 15512
rect 19628 15026 19656 15506
rect 19616 15020 19668 15026
rect 19616 14962 19668 14968
rect 19720 14346 19748 16390
rect 19800 15904 19852 15910
rect 19800 15846 19852 15852
rect 19812 15502 19840 15846
rect 19800 15496 19852 15502
rect 19800 15438 19852 15444
rect 19708 14340 19760 14346
rect 19708 14282 19760 14288
rect 19708 13932 19760 13938
rect 19760 13892 19840 13920
rect 19708 13874 19760 13880
rect 19522 13832 19578 13841
rect 19522 13767 19578 13776
rect 19524 13728 19576 13734
rect 19524 13670 19576 13676
rect 19616 13728 19668 13734
rect 19616 13670 19668 13676
rect 19536 12646 19564 13670
rect 19628 13530 19656 13670
rect 19616 13524 19668 13530
rect 19616 13466 19668 13472
rect 19708 13524 19760 13530
rect 19708 13466 19760 13472
rect 19628 13326 19656 13466
rect 19720 13326 19748 13466
rect 19616 13320 19668 13326
rect 19616 13262 19668 13268
rect 19708 13320 19760 13326
rect 19708 13262 19760 13268
rect 19812 12918 19840 13892
rect 19800 12912 19852 12918
rect 19706 12880 19762 12889
rect 19616 12844 19668 12850
rect 19800 12854 19852 12860
rect 19706 12815 19708 12824
rect 19616 12786 19668 12792
rect 19760 12815 19762 12824
rect 19708 12786 19760 12792
rect 19524 12640 19576 12646
rect 19524 12582 19576 12588
rect 19432 12436 19484 12442
rect 19432 12378 19484 12384
rect 19340 12232 19392 12238
rect 19392 12180 19564 12186
rect 19340 12174 19564 12180
rect 19352 12170 19564 12174
rect 19352 12164 19576 12170
rect 19352 12158 19524 12164
rect 19524 12106 19576 12112
rect 19340 11892 19392 11898
rect 19340 11834 19392 11840
rect 19352 11150 19380 11834
rect 19628 11694 19656 12786
rect 19904 12730 19932 16934
rect 20076 14816 20128 14822
rect 20076 14758 20128 14764
rect 19984 13728 20036 13734
rect 19984 13670 20036 13676
rect 19996 13394 20024 13670
rect 19984 13388 20036 13394
rect 19984 13330 20036 13336
rect 20088 13274 20116 14758
rect 20260 13796 20312 13802
rect 20260 13738 20312 13744
rect 19720 12702 19932 12730
rect 19996 13246 20116 13274
rect 19616 11688 19668 11694
rect 19616 11630 19668 11636
rect 19340 11144 19392 11150
rect 19340 11086 19392 11092
rect 19432 11144 19484 11150
rect 19432 11086 19484 11092
rect 19444 10130 19472 11086
rect 19616 10192 19668 10198
rect 19616 10134 19668 10140
rect 19432 10124 19484 10130
rect 19432 10066 19484 10072
rect 19628 9994 19656 10134
rect 19616 9988 19668 9994
rect 19616 9930 19668 9936
rect 19628 9382 19656 9930
rect 19616 9376 19668 9382
rect 19616 9318 19668 9324
rect 19720 8650 19748 12702
rect 19892 12640 19944 12646
rect 19892 12582 19944 12588
rect 19800 12232 19852 12238
rect 19800 12174 19852 12180
rect 19812 11354 19840 12174
rect 19800 11348 19852 11354
rect 19800 11290 19852 11296
rect 19800 11144 19852 11150
rect 19800 11086 19852 11092
rect 19812 9926 19840 11086
rect 19904 10674 19932 12582
rect 19996 11898 20024 13246
rect 20272 13190 20300 13738
rect 20364 13734 20392 17138
rect 20536 17128 20588 17134
rect 20536 17070 20588 17076
rect 20444 16720 20496 16726
rect 20444 16662 20496 16668
rect 20456 16590 20484 16662
rect 20548 16658 20576 17070
rect 20732 16658 20760 17478
rect 20824 17241 20852 17614
rect 21364 17604 21416 17610
rect 21364 17546 21416 17552
rect 20996 17536 21048 17542
rect 20996 17478 21048 17484
rect 20810 17232 20866 17241
rect 20810 17167 20812 17176
rect 20864 17167 20866 17176
rect 20904 17196 20956 17202
rect 20812 17138 20864 17144
rect 21008 17184 21036 17478
rect 20956 17156 21036 17184
rect 20904 17138 20956 17144
rect 20812 16992 20864 16998
rect 20812 16934 20864 16940
rect 20536 16652 20588 16658
rect 20536 16594 20588 16600
rect 20720 16652 20772 16658
rect 20720 16594 20772 16600
rect 20444 16584 20496 16590
rect 20444 16526 20496 16532
rect 20824 16114 20852 16934
rect 21008 16726 21036 17156
rect 20996 16720 21048 16726
rect 20996 16662 21048 16668
rect 21270 16688 21326 16697
rect 21008 16538 21036 16662
rect 21270 16623 21326 16632
rect 21008 16522 21128 16538
rect 21008 16516 21140 16522
rect 21008 16510 21088 16516
rect 21088 16458 21140 16464
rect 21284 16454 21312 16623
rect 21376 16454 21404 17546
rect 21548 17536 21600 17542
rect 21548 17478 21600 17484
rect 21560 17202 21588 17478
rect 21822 17368 21878 17377
rect 21928 17338 21956 18158
rect 22192 17808 22244 17814
rect 22192 17750 22244 17756
rect 21822 17303 21878 17312
rect 21916 17332 21968 17338
rect 21836 17202 21864 17303
rect 21916 17274 21968 17280
rect 21548 17196 21600 17202
rect 21548 17138 21600 17144
rect 21824 17196 21876 17202
rect 22100 17196 22152 17202
rect 21824 17138 21876 17144
rect 22020 17156 22100 17184
rect 21456 16992 21508 16998
rect 21456 16934 21508 16940
rect 21468 16658 21496 16934
rect 21456 16652 21508 16658
rect 21456 16594 21508 16600
rect 21640 16516 21692 16522
rect 21640 16458 21692 16464
rect 20996 16448 21048 16454
rect 20996 16390 21048 16396
rect 21272 16448 21324 16454
rect 21272 16390 21324 16396
rect 21364 16448 21416 16454
rect 21364 16390 21416 16396
rect 20536 16108 20588 16114
rect 20536 16050 20588 16056
rect 20812 16108 20864 16114
rect 20812 16050 20864 16056
rect 20548 15337 20576 16050
rect 21008 16046 21036 16390
rect 21284 16114 21312 16390
rect 21652 16114 21680 16458
rect 22020 16250 22048 17156
rect 22100 17138 22152 17144
rect 22100 16788 22152 16794
rect 22100 16730 22152 16736
rect 22112 16590 22140 16730
rect 22100 16584 22152 16590
rect 22100 16526 22152 16532
rect 22008 16244 22060 16250
rect 22008 16186 22060 16192
rect 21272 16108 21324 16114
rect 21272 16050 21324 16056
rect 21640 16108 21692 16114
rect 21640 16050 21692 16056
rect 20996 16040 21048 16046
rect 20996 15982 21048 15988
rect 21008 15570 21036 15982
rect 21088 15904 21140 15910
rect 21088 15846 21140 15852
rect 21100 15706 21128 15846
rect 21284 15706 21312 16050
rect 21364 15904 21416 15910
rect 21364 15846 21416 15852
rect 21088 15700 21140 15706
rect 21088 15642 21140 15648
rect 21272 15700 21324 15706
rect 21272 15642 21324 15648
rect 21376 15638 21404 15846
rect 21364 15632 21416 15638
rect 21364 15574 21416 15580
rect 20996 15564 21048 15570
rect 20996 15506 21048 15512
rect 21652 15502 21680 16050
rect 22112 16046 22140 16526
rect 22204 16182 22232 17750
rect 22192 16176 22244 16182
rect 22192 16118 22244 16124
rect 22100 16040 22152 16046
rect 22100 15982 22152 15988
rect 22296 15858 22324 19672
rect 22112 15830 22324 15858
rect 22112 15586 22140 15830
rect 22388 15722 22416 19722
rect 22572 19514 22600 19790
rect 22560 19508 22612 19514
rect 22560 19450 22612 19456
rect 22466 19408 22522 19417
rect 22466 19343 22468 19352
rect 22520 19343 22522 19352
rect 22468 19314 22520 19320
rect 22480 18426 22508 19314
rect 22468 18420 22520 18426
rect 22468 18362 22520 18368
rect 22572 16574 22600 19450
rect 22664 19378 22692 19858
rect 22652 19372 22704 19378
rect 22652 19314 22704 19320
rect 22756 19258 22784 20295
rect 22848 19922 22876 20470
rect 22836 19916 22888 19922
rect 22836 19858 22888 19864
rect 22020 15558 22140 15586
rect 22204 15694 22416 15722
rect 22480 16546 22600 16574
rect 22664 19230 22784 19258
rect 20720 15496 20772 15502
rect 20720 15438 20772 15444
rect 21272 15496 21324 15502
rect 21272 15438 21324 15444
rect 21456 15496 21508 15502
rect 21456 15438 21508 15444
rect 21640 15496 21692 15502
rect 21640 15438 21692 15444
rect 20534 15328 20590 15337
rect 20534 15263 20590 15272
rect 20732 15162 20760 15438
rect 20720 15156 20772 15162
rect 20720 15098 20772 15104
rect 21284 15026 21312 15438
rect 21272 15020 21324 15026
rect 21272 14962 21324 14968
rect 21468 14958 21496 15438
rect 22020 15094 22048 15558
rect 22100 15496 22152 15502
rect 22100 15438 22152 15444
rect 22008 15088 22060 15094
rect 22008 15030 22060 15036
rect 21456 14952 21508 14958
rect 21456 14894 21508 14900
rect 21824 14952 21876 14958
rect 21824 14894 21876 14900
rect 20720 14476 20772 14482
rect 20720 14418 20772 14424
rect 20628 14340 20680 14346
rect 20628 14282 20680 14288
rect 20444 14272 20496 14278
rect 20444 14214 20496 14220
rect 20536 14272 20588 14278
rect 20536 14214 20588 14220
rect 20456 13870 20484 14214
rect 20548 14074 20576 14214
rect 20536 14068 20588 14074
rect 20536 14010 20588 14016
rect 20640 13954 20668 14282
rect 20732 14074 20760 14418
rect 20720 14068 20772 14074
rect 20720 14010 20772 14016
rect 21548 14068 21600 14074
rect 21548 14010 21600 14016
rect 20548 13926 20668 13954
rect 21364 14000 21416 14006
rect 21364 13942 21416 13948
rect 20904 13932 20956 13938
rect 20548 13870 20576 13926
rect 20904 13874 20956 13880
rect 20444 13864 20496 13870
rect 20444 13806 20496 13812
rect 20536 13864 20588 13870
rect 20628 13864 20680 13870
rect 20536 13806 20588 13812
rect 20626 13832 20628 13841
rect 20916 13841 20944 13874
rect 20680 13832 20682 13841
rect 20352 13728 20404 13734
rect 20352 13670 20404 13676
rect 20352 13524 20404 13530
rect 20352 13466 20404 13472
rect 20260 13184 20312 13190
rect 20260 13126 20312 13132
rect 20168 12980 20220 12986
rect 20168 12922 20220 12928
rect 20076 12912 20128 12918
rect 20076 12854 20128 12860
rect 19984 11892 20036 11898
rect 19984 11834 20036 11840
rect 20088 11665 20116 12854
rect 20180 12764 20208 12922
rect 20364 12850 20392 13466
rect 20352 12844 20404 12850
rect 20352 12786 20404 12792
rect 20260 12776 20312 12782
rect 20180 12736 20260 12764
rect 20180 12646 20208 12736
rect 20260 12718 20312 12724
rect 20168 12640 20220 12646
rect 20168 12582 20220 12588
rect 20168 11892 20220 11898
rect 20168 11834 20220 11840
rect 20074 11656 20130 11665
rect 20074 11591 20130 11600
rect 19984 11552 20036 11558
rect 19984 11494 20036 11500
rect 19996 11354 20024 11494
rect 19984 11348 20036 11354
rect 19984 11290 20036 11296
rect 20180 11286 20208 11834
rect 20168 11280 20220 11286
rect 20168 11222 20220 11228
rect 20456 11150 20484 13806
rect 20626 13767 20682 13776
rect 20902 13832 20958 13841
rect 20902 13767 20958 13776
rect 21376 13530 21404 13942
rect 21364 13524 21416 13530
rect 21364 13466 21416 13472
rect 21180 13388 21232 13394
rect 21180 13330 21232 13336
rect 21192 12850 21220 13330
rect 21364 13252 21416 13258
rect 21364 13194 21416 13200
rect 20536 12844 20588 12850
rect 20536 12786 20588 12792
rect 20812 12844 20864 12850
rect 20996 12844 21048 12850
rect 20864 12804 20996 12832
rect 20812 12786 20864 12792
rect 20996 12786 21048 12792
rect 21180 12844 21232 12850
rect 21180 12786 21232 12792
rect 20548 12102 20576 12786
rect 20720 12640 20772 12646
rect 20720 12582 20772 12588
rect 21088 12640 21140 12646
rect 21088 12582 21140 12588
rect 20732 12306 20760 12582
rect 20720 12300 20772 12306
rect 20720 12242 20772 12248
rect 20536 12096 20588 12102
rect 20536 12038 20588 12044
rect 20444 11144 20496 11150
rect 20444 11086 20496 11092
rect 19892 10668 19944 10674
rect 19892 10610 19944 10616
rect 20260 10464 20312 10470
rect 20260 10406 20312 10412
rect 20272 10130 20300 10406
rect 20260 10124 20312 10130
rect 20260 10066 20312 10072
rect 20548 10062 20576 12038
rect 20732 11558 20760 12242
rect 21100 12238 21128 12582
rect 21376 12434 21404 13194
rect 21376 12406 21496 12434
rect 21088 12232 21140 12238
rect 21088 12174 21140 12180
rect 21100 11762 21128 12174
rect 21272 12164 21324 12170
rect 21272 12106 21324 12112
rect 21088 11756 21140 11762
rect 21088 11698 21140 11704
rect 20812 11688 20864 11694
rect 20812 11630 20864 11636
rect 20720 11552 20772 11558
rect 20720 11494 20772 11500
rect 20824 11082 20852 11630
rect 21180 11348 21232 11354
rect 21180 11290 21232 11296
rect 20812 11076 20864 11082
rect 20812 11018 20864 11024
rect 20720 11008 20772 11014
rect 20720 10950 20772 10956
rect 20732 10674 20760 10950
rect 20720 10668 20772 10674
rect 20720 10610 20772 10616
rect 20168 10056 20220 10062
rect 20168 9998 20220 10004
rect 20352 10056 20404 10062
rect 20352 9998 20404 10004
rect 20536 10056 20588 10062
rect 20536 9998 20588 10004
rect 19800 9920 19852 9926
rect 19800 9862 19852 9868
rect 19628 8622 19748 8650
rect 19432 8356 19484 8362
rect 19432 8298 19484 8304
rect 19444 7818 19472 8298
rect 19524 8288 19576 8294
rect 19628 8265 19656 8622
rect 19708 8356 19760 8362
rect 19708 8298 19760 8304
rect 19524 8230 19576 8236
rect 19614 8256 19670 8265
rect 19536 8106 19564 8230
rect 19614 8191 19670 8200
rect 19536 8078 19656 8106
rect 19628 7886 19656 8078
rect 19720 7954 19748 8298
rect 19708 7948 19760 7954
rect 19708 7890 19760 7896
rect 19524 7880 19576 7886
rect 19522 7848 19524 7857
rect 19616 7880 19668 7886
rect 19576 7848 19578 7857
rect 19156 7812 19208 7818
rect 19156 7754 19208 7760
rect 19432 7812 19484 7818
rect 19616 7822 19668 7828
rect 19522 7783 19578 7792
rect 19432 7754 19484 7760
rect 19064 7744 19116 7750
rect 19064 7686 19116 7692
rect 19248 7744 19300 7750
rect 19248 7686 19300 7692
rect 19076 7410 19104 7686
rect 19064 7404 19116 7410
rect 19064 7346 19116 7352
rect 19260 7342 19288 7686
rect 19812 7342 19840 9862
rect 20180 9586 20208 9998
rect 20168 9580 20220 9586
rect 20168 9522 20220 9528
rect 19984 9376 20036 9382
rect 19984 9318 20036 9324
rect 19996 8566 20024 9318
rect 19984 8560 20036 8566
rect 19984 8502 20036 8508
rect 20180 8362 20208 9522
rect 20260 8424 20312 8430
rect 20260 8366 20312 8372
rect 20168 8356 20220 8362
rect 20168 8298 20220 8304
rect 19892 8288 19944 8294
rect 20272 8242 20300 8366
rect 19892 8230 19944 8236
rect 19904 8090 19932 8230
rect 19996 8214 20300 8242
rect 19892 8084 19944 8090
rect 19892 8026 19944 8032
rect 19996 7886 20024 8214
rect 20074 8120 20130 8129
rect 20074 8055 20076 8064
rect 20128 8055 20130 8064
rect 20076 8026 20128 8032
rect 19984 7880 20036 7886
rect 19984 7822 20036 7828
rect 20074 7576 20130 7585
rect 20074 7511 20076 7520
rect 20128 7511 20130 7520
rect 20076 7482 20128 7488
rect 19248 7336 19300 7342
rect 19248 7278 19300 7284
rect 19800 7336 19852 7342
rect 19800 7278 19852 7284
rect 20364 6866 20392 9998
rect 20824 9994 20852 11018
rect 21192 10674 21220 11290
rect 21284 11150 21312 12106
rect 21364 11348 21416 11354
rect 21364 11290 21416 11296
rect 21376 11150 21404 11290
rect 21272 11144 21324 11150
rect 21272 11086 21324 11092
rect 21364 11144 21416 11150
rect 21364 11086 21416 11092
rect 21180 10668 21232 10674
rect 21180 10610 21232 10616
rect 20904 10532 20956 10538
rect 20904 10474 20956 10480
rect 20812 9988 20864 9994
rect 20812 9930 20864 9936
rect 20720 9920 20772 9926
rect 20720 9862 20772 9868
rect 20732 9382 20760 9862
rect 20824 9654 20852 9930
rect 20812 9648 20864 9654
rect 20812 9590 20864 9596
rect 20916 9466 20944 10474
rect 20824 9438 20944 9466
rect 20720 9376 20772 9382
rect 20720 9318 20772 9324
rect 20628 8288 20680 8294
rect 20628 8230 20680 8236
rect 20640 7886 20668 8230
rect 20444 7880 20496 7886
rect 20444 7822 20496 7828
rect 20536 7880 20588 7886
rect 20536 7822 20588 7828
rect 20628 7880 20680 7886
rect 20628 7822 20680 7828
rect 20456 7274 20484 7822
rect 20548 7546 20576 7822
rect 20536 7540 20588 7546
rect 20536 7482 20588 7488
rect 20548 7342 20576 7482
rect 20824 7410 20852 9438
rect 21088 9376 21140 9382
rect 21088 9318 21140 9324
rect 20904 8492 20956 8498
rect 20904 8434 20956 8440
rect 20916 7449 20944 8434
rect 20996 8288 21048 8294
rect 20996 8230 21048 8236
rect 21008 7993 21036 8230
rect 20994 7984 21050 7993
rect 20994 7919 21050 7928
rect 20902 7440 20958 7449
rect 20812 7404 20864 7410
rect 20902 7375 20904 7384
rect 20812 7346 20864 7352
rect 20956 7375 20958 7384
rect 21008 7392 21036 7919
rect 21100 7886 21128 9318
rect 21192 8294 21220 10610
rect 21376 9674 21404 11086
rect 21468 9994 21496 12406
rect 21560 11354 21588 14010
rect 21640 13932 21692 13938
rect 21640 13874 21692 13880
rect 21652 13530 21680 13874
rect 21640 13524 21692 13530
rect 21640 13466 21692 13472
rect 21732 13524 21784 13530
rect 21732 13466 21784 13472
rect 21640 13184 21692 13190
rect 21640 13126 21692 13132
rect 21652 12918 21680 13126
rect 21640 12912 21692 12918
rect 21640 12854 21692 12860
rect 21548 11348 21600 11354
rect 21548 11290 21600 11296
rect 21548 11212 21600 11218
rect 21548 11154 21600 11160
rect 21560 10674 21588 11154
rect 21744 10742 21772 13466
rect 21836 13462 21864 14894
rect 21824 13456 21876 13462
rect 21824 13398 21876 13404
rect 21836 12889 21864 13398
rect 22112 13326 22140 15438
rect 22204 13530 22232 15694
rect 22376 15632 22428 15638
rect 22376 15574 22428 15580
rect 22388 14906 22416 15574
rect 22296 14878 22416 14906
rect 22296 14521 22324 14878
rect 22282 14512 22338 14521
rect 22282 14447 22338 14456
rect 22376 14476 22428 14482
rect 22296 13938 22324 14447
rect 22376 14418 22428 14424
rect 22388 14006 22416 14418
rect 22376 14000 22428 14006
rect 22376 13942 22428 13948
rect 22284 13932 22336 13938
rect 22284 13874 22336 13880
rect 22282 13832 22338 13841
rect 22282 13767 22338 13776
rect 22192 13524 22244 13530
rect 22192 13466 22244 13472
rect 22100 13320 22152 13326
rect 22100 13262 22152 13268
rect 22192 13320 22244 13326
rect 22192 13262 22244 13268
rect 21916 13252 21968 13258
rect 21916 13194 21968 13200
rect 21822 12880 21878 12889
rect 21822 12815 21878 12824
rect 21928 12832 21956 13194
rect 22008 12844 22060 12850
rect 21928 12804 22008 12832
rect 22008 12786 22060 12792
rect 21732 10736 21784 10742
rect 21732 10678 21784 10684
rect 21548 10668 21600 10674
rect 21548 10610 21600 10616
rect 21744 10538 21772 10678
rect 21824 10600 21876 10606
rect 21824 10542 21876 10548
rect 21916 10600 21968 10606
rect 21916 10542 21968 10548
rect 21732 10532 21784 10538
rect 21732 10474 21784 10480
rect 21456 9988 21508 9994
rect 21456 9930 21508 9936
rect 21468 9722 21496 9930
rect 21836 9722 21864 10542
rect 21284 9646 21404 9674
rect 21456 9716 21508 9722
rect 21456 9658 21508 9664
rect 21824 9716 21876 9722
rect 21824 9658 21876 9664
rect 21180 8288 21232 8294
rect 21180 8230 21232 8236
rect 21284 8022 21312 9646
rect 21272 8016 21324 8022
rect 21272 7958 21324 7964
rect 21180 7948 21232 7954
rect 21180 7890 21232 7896
rect 21088 7880 21140 7886
rect 21088 7822 21140 7828
rect 21192 7478 21220 7890
rect 21180 7472 21232 7478
rect 21180 7414 21232 7420
rect 21088 7404 21140 7410
rect 21008 7364 21088 7392
rect 20904 7346 20956 7352
rect 21088 7346 21140 7352
rect 20536 7336 20588 7342
rect 20536 7278 20588 7284
rect 20444 7268 20496 7274
rect 20444 7210 20496 7216
rect 21180 7200 21232 7206
rect 21284 7188 21312 7958
rect 21232 7160 21312 7188
rect 21364 7200 21416 7206
rect 21180 7142 21232 7148
rect 21364 7142 21416 7148
rect 21376 7002 21404 7142
rect 21364 6996 21416 7002
rect 21364 6938 21416 6944
rect 18972 6860 19024 6866
rect 18972 6802 19024 6808
rect 20352 6860 20404 6866
rect 20352 6802 20404 6808
rect 21468 6798 21496 9658
rect 21928 9330 21956 10542
rect 22020 9450 22048 12786
rect 22112 12782 22140 13262
rect 22100 12776 22152 12782
rect 22100 12718 22152 12724
rect 22204 12714 22232 13262
rect 22296 13258 22324 13767
rect 22284 13252 22336 13258
rect 22284 13194 22336 13200
rect 22296 12918 22324 13194
rect 22388 12986 22416 13942
rect 22480 13938 22508 16546
rect 22560 16108 22612 16114
rect 22560 16050 22612 16056
rect 22572 13938 22600 16050
rect 22664 15638 22692 19230
rect 22848 18834 22876 19858
rect 22940 19854 22968 21422
rect 23020 21344 23072 21350
rect 23020 21286 23072 21292
rect 23032 20942 23060 21286
rect 23020 20936 23072 20942
rect 23020 20878 23072 20884
rect 22928 19848 22980 19854
rect 22928 19790 22980 19796
rect 23020 19372 23072 19378
rect 22940 19320 23020 19334
rect 22940 19314 23072 19320
rect 22940 19306 23060 19314
rect 22836 18828 22888 18834
rect 22836 18770 22888 18776
rect 22744 18420 22796 18426
rect 22744 18362 22796 18368
rect 22756 16114 22784 18362
rect 22848 18290 22876 18770
rect 22836 18284 22888 18290
rect 22836 18226 22888 18232
rect 22940 17746 22968 19306
rect 23124 17746 23152 21490
rect 23308 20942 23336 21626
rect 23938 21312 23994 21321
rect 23938 21247 23994 21256
rect 23952 21146 23980 21247
rect 23940 21140 23992 21146
rect 23940 21082 23992 21088
rect 23296 20936 23348 20942
rect 23296 20878 23348 20884
rect 23388 20936 23440 20942
rect 23388 20878 23440 20884
rect 23400 20058 23428 20878
rect 23572 20868 23624 20874
rect 23572 20810 23624 20816
rect 23388 20052 23440 20058
rect 23388 19994 23440 20000
rect 23296 19984 23348 19990
rect 23348 19932 23428 19938
rect 23296 19926 23428 19932
rect 23308 19910 23428 19926
rect 23296 19848 23348 19854
rect 23296 19790 23348 19796
rect 23308 19378 23336 19790
rect 23400 19378 23428 19910
rect 23584 19514 23612 20810
rect 23756 20256 23808 20262
rect 23756 20198 23808 20204
rect 23664 19780 23716 19786
rect 23664 19722 23716 19728
rect 23572 19508 23624 19514
rect 23572 19450 23624 19456
rect 23676 19446 23704 19722
rect 23664 19440 23716 19446
rect 23664 19382 23716 19388
rect 23296 19372 23348 19378
rect 23296 19314 23348 19320
rect 23388 19372 23440 19378
rect 23388 19314 23440 19320
rect 23400 17898 23428 19314
rect 23480 19168 23532 19174
rect 23480 19110 23532 19116
rect 23216 17870 23428 17898
rect 22928 17740 22980 17746
rect 22928 17682 22980 17688
rect 23112 17740 23164 17746
rect 23112 17682 23164 17688
rect 22940 17066 22968 17682
rect 23216 17678 23244 17870
rect 23296 17740 23348 17746
rect 23296 17682 23348 17688
rect 23204 17672 23256 17678
rect 23204 17614 23256 17620
rect 23216 17542 23244 17614
rect 23204 17536 23256 17542
rect 23204 17478 23256 17484
rect 23204 17196 23256 17202
rect 23204 17138 23256 17144
rect 22928 17060 22980 17066
rect 22928 17002 22980 17008
rect 22744 16108 22796 16114
rect 22744 16050 22796 16056
rect 22928 16108 22980 16114
rect 22928 16050 22980 16056
rect 22652 15632 22704 15638
rect 22652 15574 22704 15580
rect 22756 14770 22784 16050
rect 22940 15638 22968 16050
rect 22928 15632 22980 15638
rect 22928 15574 22980 15580
rect 23216 15502 23244 17138
rect 23308 15994 23336 17682
rect 23492 17202 23520 19110
rect 23480 17196 23532 17202
rect 23480 17138 23532 17144
rect 23676 17134 23704 19382
rect 23768 18358 23796 20198
rect 23952 19258 23980 21082
rect 24412 20942 24440 23122
rect 24688 22030 24716 24142
rect 24780 24138 24808 24754
rect 24872 24750 24900 26318
rect 24964 25430 24992 26454
rect 25320 26376 25372 26382
rect 25320 26318 25372 26324
rect 25412 26376 25464 26382
rect 25516 26364 25544 27406
rect 25780 27328 25832 27334
rect 25780 27270 25832 27276
rect 25596 26852 25648 26858
rect 25596 26794 25648 26800
rect 25464 26336 25544 26364
rect 25412 26318 25464 26324
rect 25136 26240 25188 26246
rect 25136 26182 25188 26188
rect 24952 25424 25004 25430
rect 24952 25366 25004 25372
rect 24964 24886 24992 25366
rect 24952 24880 25004 24886
rect 24952 24822 25004 24828
rect 25148 24750 25176 26182
rect 24860 24744 24912 24750
rect 24860 24686 24912 24692
rect 24952 24744 25004 24750
rect 24952 24686 25004 24692
rect 25136 24744 25188 24750
rect 25136 24686 25188 24692
rect 24964 24410 24992 24686
rect 24952 24404 25004 24410
rect 24952 24346 25004 24352
rect 24952 24268 25004 24274
rect 24952 24210 25004 24216
rect 24768 24132 24820 24138
rect 24768 24074 24820 24080
rect 24964 23866 24992 24210
rect 25332 24138 25360 26318
rect 25320 24132 25372 24138
rect 25320 24074 25372 24080
rect 24952 23860 25004 23866
rect 24952 23802 25004 23808
rect 25332 23798 25360 24074
rect 25136 23792 25188 23798
rect 25136 23734 25188 23740
rect 25320 23792 25372 23798
rect 25320 23734 25372 23740
rect 25044 23656 25096 23662
rect 25044 23598 25096 23604
rect 24676 22024 24728 22030
rect 24676 21966 24728 21972
rect 25056 21978 25084 23598
rect 25148 23050 25176 23734
rect 25136 23044 25188 23050
rect 25136 22986 25188 22992
rect 25148 22953 25176 22986
rect 25134 22944 25190 22953
rect 25134 22879 25190 22888
rect 25424 22438 25452 26318
rect 25504 25696 25556 25702
rect 25504 25638 25556 25644
rect 25516 24274 25544 25638
rect 25608 24614 25636 26794
rect 25792 26382 25820 27270
rect 25884 27130 25912 28494
rect 25964 27668 26016 27674
rect 25964 27610 26016 27616
rect 25976 27470 26004 27610
rect 25964 27464 26016 27470
rect 25964 27406 26016 27412
rect 25964 27328 26016 27334
rect 25964 27270 26016 27276
rect 25872 27124 25924 27130
rect 25872 27066 25924 27072
rect 25870 27024 25926 27033
rect 25976 26994 26004 27270
rect 26068 27130 26096 28494
rect 26148 28484 26200 28490
rect 26148 28426 26200 28432
rect 26056 27124 26108 27130
rect 26056 27066 26108 27072
rect 25870 26959 25872 26968
rect 25924 26959 25926 26968
rect 25964 26988 26016 26994
rect 25872 26930 25924 26936
rect 25964 26930 26016 26936
rect 26160 26858 26188 28426
rect 26240 27940 26292 27946
rect 26240 27882 26292 27888
rect 26252 27402 26280 27882
rect 26804 27674 26832 28494
rect 27160 28076 27212 28082
rect 27160 28018 27212 28024
rect 27172 27674 27200 28018
rect 28000 27946 28028 30790
rect 28354 30676 28410 30790
rect 28736 30790 29054 30818
rect 28736 28218 28764 30790
rect 28998 30676 29054 30790
rect 28724 28212 28776 28218
rect 28724 28154 28776 28160
rect 27988 27940 28040 27946
rect 27988 27882 28040 27888
rect 26792 27668 26844 27674
rect 26792 27610 26844 27616
rect 27160 27668 27212 27674
rect 27160 27610 27212 27616
rect 26330 27568 26386 27577
rect 26330 27503 26332 27512
rect 26384 27503 26386 27512
rect 26332 27474 26384 27480
rect 26240 27396 26292 27402
rect 26240 27338 26292 27344
rect 26252 26994 26280 27338
rect 26240 26988 26292 26994
rect 26240 26930 26292 26936
rect 26148 26852 26200 26858
rect 26148 26794 26200 26800
rect 26252 26586 26280 26930
rect 26240 26580 26292 26586
rect 26240 26522 26292 26528
rect 26344 26432 26372 27474
rect 26792 27464 26844 27470
rect 26792 27406 26844 27412
rect 26804 27062 26832 27406
rect 26792 27056 26844 27062
rect 26792 26998 26844 27004
rect 26804 26586 26832 26998
rect 26792 26580 26844 26586
rect 26792 26522 26844 26528
rect 27712 26512 27764 26518
rect 27712 26454 27764 26460
rect 26160 26404 26372 26432
rect 25780 26376 25832 26382
rect 25832 26336 26004 26364
rect 25780 26318 25832 26324
rect 25780 26240 25832 26246
rect 25780 26182 25832 26188
rect 25792 26042 25820 26182
rect 25780 26036 25832 26042
rect 25780 25978 25832 25984
rect 25780 25900 25832 25906
rect 25780 25842 25832 25848
rect 25596 24608 25648 24614
rect 25596 24550 25648 24556
rect 25504 24268 25556 24274
rect 25504 24210 25556 24216
rect 25608 24138 25636 24550
rect 25688 24200 25740 24206
rect 25792 24188 25820 25842
rect 25872 25696 25924 25702
rect 25872 25638 25924 25644
rect 25884 25294 25912 25638
rect 25976 25362 26004 26336
rect 25964 25356 26016 25362
rect 25964 25298 26016 25304
rect 25872 25288 25924 25294
rect 26160 25276 26188 26404
rect 26700 26376 26752 26382
rect 26700 26318 26752 26324
rect 27528 26376 27580 26382
rect 27528 26318 27580 26324
rect 26240 26308 26292 26314
rect 26240 26250 26292 26256
rect 26332 26308 26384 26314
rect 26332 26250 26384 26256
rect 26252 25974 26280 26250
rect 26240 25968 26292 25974
rect 26240 25910 26292 25916
rect 26344 25906 26372 26250
rect 26332 25900 26384 25906
rect 26332 25842 26384 25848
rect 26240 25288 26292 25294
rect 26160 25248 26240 25276
rect 25872 25230 25924 25236
rect 26240 25230 26292 25236
rect 25872 24812 25924 24818
rect 25872 24754 25924 24760
rect 25884 24614 25912 24754
rect 26056 24744 26108 24750
rect 25976 24704 26056 24732
rect 25872 24608 25924 24614
rect 25872 24550 25924 24556
rect 25884 24342 25912 24550
rect 25872 24336 25924 24342
rect 25872 24278 25924 24284
rect 25872 24200 25924 24206
rect 25792 24160 25872 24188
rect 25688 24142 25740 24148
rect 25872 24142 25924 24148
rect 25504 24132 25556 24138
rect 25504 24074 25556 24080
rect 25596 24132 25648 24138
rect 25596 24074 25648 24080
rect 25516 23662 25544 24074
rect 25596 23724 25648 23730
rect 25700 23712 25728 24142
rect 25884 23866 25912 24142
rect 25976 24120 26004 24704
rect 26056 24686 26108 24692
rect 26148 24200 26200 24206
rect 26148 24142 26200 24148
rect 26056 24132 26108 24138
rect 25976 24092 26056 24120
rect 25872 23860 25924 23866
rect 25872 23802 25924 23808
rect 25648 23684 25728 23712
rect 25596 23666 25648 23672
rect 25504 23656 25556 23662
rect 25504 23598 25556 23604
rect 25700 23338 25728 23684
rect 25608 23310 25728 23338
rect 25504 22976 25556 22982
rect 25504 22918 25556 22924
rect 25412 22432 25464 22438
rect 25412 22374 25464 22380
rect 25320 22024 25372 22030
rect 25056 21950 25176 21978
rect 25320 21966 25372 21972
rect 25044 21888 25096 21894
rect 25044 21830 25096 21836
rect 24952 21684 25004 21690
rect 24952 21626 25004 21632
rect 24964 21554 24992 21626
rect 24952 21548 25004 21554
rect 24952 21490 25004 21496
rect 25056 21146 25084 21830
rect 25148 21486 25176 21950
rect 25136 21480 25188 21486
rect 25136 21422 25188 21428
rect 25148 21350 25176 21422
rect 25332 21418 25360 21966
rect 25424 21622 25452 22374
rect 25516 21962 25544 22918
rect 25504 21956 25556 21962
rect 25504 21898 25556 21904
rect 25412 21616 25464 21622
rect 25412 21558 25464 21564
rect 25320 21412 25372 21418
rect 25320 21354 25372 21360
rect 25136 21344 25188 21350
rect 25516 21298 25544 21898
rect 25608 21894 25636 23310
rect 25976 22982 26004 24092
rect 26056 24074 26108 24080
rect 26160 23118 26188 24142
rect 26252 23254 26280 25230
rect 26344 24410 26372 25842
rect 26712 25702 26740 26318
rect 27540 26042 27568 26318
rect 27528 26036 27580 26042
rect 27528 25978 27580 25984
rect 27160 25968 27212 25974
rect 27724 25945 27752 26454
rect 27160 25910 27212 25916
rect 27710 25936 27766 25945
rect 26976 25764 27028 25770
rect 26976 25706 27028 25712
rect 26424 25696 26476 25702
rect 26424 25638 26476 25644
rect 26700 25696 26752 25702
rect 26700 25638 26752 25644
rect 26436 25226 26464 25638
rect 26424 25220 26476 25226
rect 26424 25162 26476 25168
rect 26516 25152 26568 25158
rect 26516 25094 26568 25100
rect 26528 24750 26556 25094
rect 26792 24880 26844 24886
rect 26792 24822 26844 24828
rect 26516 24744 26568 24750
rect 26516 24686 26568 24692
rect 26332 24404 26384 24410
rect 26332 24346 26384 24352
rect 26528 24206 26556 24686
rect 26516 24200 26568 24206
rect 26516 24142 26568 24148
rect 26240 23248 26292 23254
rect 26240 23190 26292 23196
rect 26148 23112 26200 23118
rect 26148 23054 26200 23060
rect 25964 22976 26016 22982
rect 25964 22918 26016 22924
rect 25976 22642 26004 22918
rect 26160 22642 26188 23054
rect 25688 22636 25740 22642
rect 25688 22578 25740 22584
rect 25964 22636 26016 22642
rect 25964 22578 26016 22584
rect 26148 22636 26200 22642
rect 26148 22578 26200 22584
rect 25700 22030 25728 22578
rect 26252 22438 26280 23190
rect 26424 22772 26476 22778
rect 26424 22714 26476 22720
rect 25964 22432 26016 22438
rect 25964 22374 26016 22380
rect 26240 22432 26292 22438
rect 26240 22374 26292 22380
rect 25780 22092 25832 22098
rect 25780 22034 25832 22040
rect 25688 22024 25740 22030
rect 25688 21966 25740 21972
rect 25792 21894 25820 22034
rect 25596 21888 25648 21894
rect 25596 21830 25648 21836
rect 25780 21888 25832 21894
rect 25780 21830 25832 21836
rect 25608 21486 25636 21830
rect 25688 21548 25740 21554
rect 25688 21490 25740 21496
rect 25596 21480 25648 21486
rect 25596 21422 25648 21428
rect 25700 21298 25728 21490
rect 25792 21468 25820 21830
rect 25976 21690 26004 22374
rect 26252 22234 26280 22374
rect 26240 22228 26292 22234
rect 26240 22170 26292 22176
rect 26148 22160 26200 22166
rect 26148 22102 26200 22108
rect 26056 21956 26108 21962
rect 26056 21898 26108 21904
rect 25964 21684 26016 21690
rect 25964 21626 26016 21632
rect 25792 21440 25912 21468
rect 25136 21286 25188 21292
rect 25044 21140 25096 21146
rect 25044 21082 25096 21088
rect 24308 20936 24360 20942
rect 24308 20878 24360 20884
rect 24400 20936 24452 20942
rect 24400 20878 24452 20884
rect 24216 20800 24268 20806
rect 24216 20742 24268 20748
rect 24228 20602 24256 20742
rect 24216 20596 24268 20602
rect 24216 20538 24268 20544
rect 24032 20256 24084 20262
rect 24032 20198 24084 20204
rect 24044 19786 24072 20198
rect 24032 19780 24084 19786
rect 24032 19722 24084 19728
rect 24044 19378 24072 19722
rect 24124 19712 24176 19718
rect 24124 19654 24176 19660
rect 24032 19372 24084 19378
rect 24032 19314 24084 19320
rect 23952 19230 24072 19258
rect 23756 18352 23808 18358
rect 23756 18294 23808 18300
rect 23768 18086 23796 18294
rect 23756 18080 23808 18086
rect 23756 18022 23808 18028
rect 23848 17672 23900 17678
rect 23848 17614 23900 17620
rect 23756 17604 23808 17610
rect 23756 17546 23808 17552
rect 23768 17202 23796 17546
rect 23756 17196 23808 17202
rect 23756 17138 23808 17144
rect 23664 17128 23716 17134
rect 23664 17070 23716 17076
rect 23388 16448 23440 16454
rect 23388 16390 23440 16396
rect 23400 16182 23428 16390
rect 23388 16176 23440 16182
rect 23388 16118 23440 16124
rect 23860 16114 23888 17614
rect 23940 17128 23992 17134
rect 23940 17070 23992 17076
rect 23572 16108 23624 16114
rect 23572 16050 23624 16056
rect 23848 16108 23900 16114
rect 23848 16050 23900 16056
rect 23388 16040 23440 16046
rect 23308 15988 23388 15994
rect 23308 15982 23440 15988
rect 23308 15966 23428 15982
rect 23204 15496 23256 15502
rect 23204 15438 23256 15444
rect 22664 14742 22784 14770
rect 23020 14816 23072 14822
rect 23020 14758 23072 14764
rect 22468 13932 22520 13938
rect 22468 13874 22520 13880
rect 22560 13932 22612 13938
rect 22560 13874 22612 13880
rect 22560 13796 22612 13802
rect 22560 13738 22612 13744
rect 22572 13258 22600 13738
rect 22560 13252 22612 13258
rect 22560 13194 22612 13200
rect 22376 12980 22428 12986
rect 22376 12922 22428 12928
rect 22284 12912 22336 12918
rect 22284 12854 22336 12860
rect 22192 12708 22244 12714
rect 22192 12650 22244 12656
rect 22192 10260 22244 10266
rect 22192 10202 22244 10208
rect 22204 9586 22232 10202
rect 22296 9654 22324 12854
rect 22664 11830 22692 14742
rect 22836 14272 22888 14278
rect 22836 14214 22888 14220
rect 22744 13388 22796 13394
rect 22744 13330 22796 13336
rect 22756 12986 22784 13330
rect 22744 12980 22796 12986
rect 22744 12922 22796 12928
rect 22848 12918 22876 14214
rect 23032 13938 23060 14758
rect 23296 14340 23348 14346
rect 23296 14282 23348 14288
rect 23020 13932 23072 13938
rect 23020 13874 23072 13880
rect 22928 13796 22980 13802
rect 22928 13738 22980 13744
rect 22940 13394 22968 13738
rect 23308 13530 23336 14282
rect 23400 14074 23428 15966
rect 23584 15706 23612 16050
rect 23572 15700 23624 15706
rect 23572 15642 23624 15648
rect 23756 15496 23808 15502
rect 23756 15438 23808 15444
rect 23768 14550 23796 15438
rect 23756 14544 23808 14550
rect 23756 14486 23808 14492
rect 23860 14278 23888 16050
rect 23848 14272 23900 14278
rect 23848 14214 23900 14220
rect 23388 14068 23440 14074
rect 23388 14010 23440 14016
rect 23480 13932 23532 13938
rect 23480 13874 23532 13880
rect 23388 13728 23440 13734
rect 23388 13670 23440 13676
rect 23296 13524 23348 13530
rect 23296 13466 23348 13472
rect 23400 13410 23428 13670
rect 22928 13388 22980 13394
rect 22928 13330 22980 13336
rect 23204 13388 23256 13394
rect 23204 13330 23256 13336
rect 23308 13382 23428 13410
rect 22836 12912 22888 12918
rect 22836 12854 22888 12860
rect 23216 12646 23244 13330
rect 23308 12646 23336 13382
rect 23388 12844 23440 12850
rect 23388 12786 23440 12792
rect 23204 12640 23256 12646
rect 23204 12582 23256 12588
rect 23296 12640 23348 12646
rect 23296 12582 23348 12588
rect 22652 11824 22704 11830
rect 22652 11766 22704 11772
rect 23204 11144 23256 11150
rect 23204 11086 23256 11092
rect 23216 10470 23244 11086
rect 23204 10464 23256 10470
rect 23204 10406 23256 10412
rect 22284 9648 22336 9654
rect 22284 9590 22336 9596
rect 22558 9616 22614 9625
rect 22192 9580 22244 9586
rect 22192 9522 22244 9528
rect 22008 9444 22060 9450
rect 22008 9386 22060 9392
rect 21928 9302 22048 9330
rect 22020 8430 22048 9302
rect 22008 8424 22060 8430
rect 22008 8366 22060 8372
rect 21548 7880 21600 7886
rect 21548 7822 21600 7828
rect 21560 7002 21588 7822
rect 21640 7812 21692 7818
rect 21640 7754 21692 7760
rect 21652 7410 21680 7754
rect 21732 7744 21784 7750
rect 21732 7686 21784 7692
rect 21640 7404 21692 7410
rect 21640 7346 21692 7352
rect 21744 7342 21772 7686
rect 22020 7410 22048 8366
rect 22296 8294 22324 9590
rect 22558 9551 22560 9560
rect 22612 9551 22614 9560
rect 22560 9522 22612 9528
rect 22376 9512 22428 9518
rect 22374 9480 22376 9489
rect 22428 9480 22430 9489
rect 22374 9415 22430 9424
rect 22284 8288 22336 8294
rect 22284 8230 22336 8236
rect 22192 8084 22244 8090
rect 22192 8026 22244 8032
rect 22204 7585 22232 8026
rect 22296 7857 22324 8230
rect 22282 7848 22338 7857
rect 22282 7783 22338 7792
rect 22190 7576 22246 7585
rect 22190 7511 22246 7520
rect 22296 7410 22324 7783
rect 22008 7404 22060 7410
rect 22008 7346 22060 7352
rect 22284 7404 22336 7410
rect 22284 7346 22336 7352
rect 21732 7336 21784 7342
rect 21732 7278 21784 7284
rect 22388 7274 22416 9415
rect 23400 9178 23428 12786
rect 23492 12102 23520 13874
rect 23860 13870 23888 14214
rect 23572 13864 23624 13870
rect 23572 13806 23624 13812
rect 23848 13864 23900 13870
rect 23848 13806 23900 13812
rect 23584 13530 23612 13806
rect 23572 13524 23624 13530
rect 23572 13466 23624 13472
rect 23756 13184 23808 13190
rect 23756 13126 23808 13132
rect 23572 12776 23624 12782
rect 23572 12718 23624 12724
rect 23480 12096 23532 12102
rect 23480 12038 23532 12044
rect 23584 11898 23612 12718
rect 23572 11892 23624 11898
rect 23572 11834 23624 11840
rect 23664 11144 23716 11150
rect 23664 11086 23716 11092
rect 23676 10538 23704 11086
rect 23768 10742 23796 13126
rect 23848 11756 23900 11762
rect 23848 11698 23900 11704
rect 23860 10810 23888 11698
rect 23952 11286 23980 17070
rect 24044 15502 24072 19230
rect 24032 15496 24084 15502
rect 24030 15464 24032 15473
rect 24084 15464 24086 15473
rect 24030 15399 24086 15408
rect 24136 14346 24164 19654
rect 24216 17672 24268 17678
rect 24216 17614 24268 17620
rect 24228 17338 24256 17614
rect 24216 17332 24268 17338
rect 24216 17274 24268 17280
rect 24320 16574 24348 20878
rect 25044 20800 25096 20806
rect 25044 20742 25096 20748
rect 25056 20602 25084 20742
rect 25044 20596 25096 20602
rect 25044 20538 25096 20544
rect 24860 18624 24912 18630
rect 24860 18566 24912 18572
rect 24872 18086 24900 18566
rect 25148 18426 25176 21286
rect 25424 21270 25728 21298
rect 25780 21344 25832 21350
rect 25780 21286 25832 21292
rect 25320 20936 25372 20942
rect 25320 20878 25372 20884
rect 25228 20800 25280 20806
rect 25228 20742 25280 20748
rect 25240 18698 25268 20742
rect 25332 19922 25360 20878
rect 25320 19916 25372 19922
rect 25320 19858 25372 19864
rect 25228 18692 25280 18698
rect 25228 18634 25280 18640
rect 25136 18420 25188 18426
rect 25136 18362 25188 18368
rect 24860 18080 24912 18086
rect 24860 18022 24912 18028
rect 24492 17672 24544 17678
rect 24492 17614 24544 17620
rect 24400 17536 24452 17542
rect 24400 17478 24452 17484
rect 24412 17270 24440 17478
rect 24400 17264 24452 17270
rect 24400 17206 24452 17212
rect 24504 17202 24532 17614
rect 24872 17610 24900 18022
rect 24860 17604 24912 17610
rect 24860 17546 24912 17552
rect 24768 17536 24820 17542
rect 24768 17478 24820 17484
rect 24780 17202 24808 17478
rect 24492 17196 24544 17202
rect 24492 17138 24544 17144
rect 24768 17196 24820 17202
rect 24768 17138 24820 17144
rect 24228 16546 24348 16574
rect 24228 15502 24256 16546
rect 24504 15706 24532 17138
rect 25320 16516 25372 16522
rect 25320 16458 25372 16464
rect 24860 16448 24912 16454
rect 24860 16390 24912 16396
rect 24492 15700 24544 15706
rect 24492 15642 24544 15648
rect 24584 15700 24636 15706
rect 24584 15642 24636 15648
rect 24596 15570 24624 15642
rect 24584 15564 24636 15570
rect 24584 15506 24636 15512
rect 24216 15496 24268 15502
rect 24216 15438 24268 15444
rect 24124 14340 24176 14346
rect 24124 14282 24176 14288
rect 24032 13252 24084 13258
rect 24032 13194 24084 13200
rect 24044 12918 24072 13194
rect 24032 12912 24084 12918
rect 24032 12854 24084 12860
rect 24044 11778 24072 12854
rect 24136 12434 24164 14282
rect 24228 13326 24256 15438
rect 24596 15026 24624 15506
rect 24872 15434 24900 16390
rect 25332 16250 25360 16458
rect 25320 16244 25372 16250
rect 25320 16186 25372 16192
rect 25136 15496 25188 15502
rect 25136 15438 25188 15444
rect 24860 15428 24912 15434
rect 24860 15370 24912 15376
rect 24584 15020 24636 15026
rect 24584 14962 24636 14968
rect 24596 14414 24624 14962
rect 24860 14612 24912 14618
rect 24860 14554 24912 14560
rect 24768 14544 24820 14550
rect 24768 14486 24820 14492
rect 24584 14408 24636 14414
rect 24584 14350 24636 14356
rect 24596 14074 24624 14350
rect 24584 14068 24636 14074
rect 24584 14010 24636 14016
rect 24780 13326 24808 14486
rect 24216 13320 24268 13326
rect 24584 13320 24636 13326
rect 24216 13262 24268 13268
rect 24582 13288 24584 13297
rect 24768 13320 24820 13326
rect 24636 13288 24638 13297
rect 24768 13262 24820 13268
rect 24582 13223 24638 13232
rect 24872 12986 24900 14554
rect 25148 14482 25176 15438
rect 25424 14618 25452 21270
rect 25792 20466 25820 21286
rect 25884 20874 25912 21440
rect 26068 21146 26096 21898
rect 26160 21690 26188 22102
rect 26148 21684 26200 21690
rect 26148 21626 26200 21632
rect 26252 21622 26280 22170
rect 26436 22098 26464 22714
rect 26424 22092 26476 22098
rect 26424 22034 26476 22040
rect 26240 21616 26292 21622
rect 26240 21558 26292 21564
rect 26148 21412 26200 21418
rect 26148 21354 26200 21360
rect 26056 21140 26108 21146
rect 26056 21082 26108 21088
rect 25872 20868 25924 20874
rect 25872 20810 25924 20816
rect 25872 20596 25924 20602
rect 25872 20538 25924 20544
rect 25780 20460 25832 20466
rect 25780 20402 25832 20408
rect 25884 19786 25912 20538
rect 26160 20466 26188 21354
rect 26252 20602 26280 21558
rect 26804 21400 26832 24822
rect 26988 24818 27016 25706
rect 27172 25498 27200 25910
rect 27710 25871 27766 25880
rect 27160 25492 27212 25498
rect 27160 25434 27212 25440
rect 27710 25256 27766 25265
rect 27160 25220 27212 25226
rect 27710 25191 27766 25200
rect 27160 25162 27212 25168
rect 26976 24812 27028 24818
rect 26976 24754 27028 24760
rect 26884 24132 26936 24138
rect 26884 24074 26936 24080
rect 26896 23866 26924 24074
rect 26884 23860 26936 23866
rect 26884 23802 26936 23808
rect 26896 23050 26924 23802
rect 26884 23044 26936 23050
rect 26884 22986 26936 22992
rect 26896 22710 26924 22986
rect 26884 22704 26936 22710
rect 26884 22646 26936 22652
rect 26988 21894 27016 24754
rect 27172 24614 27200 25162
rect 27724 25158 27752 25191
rect 27712 25152 27764 25158
rect 27712 25094 27764 25100
rect 27160 24608 27212 24614
rect 27712 24608 27764 24614
rect 27160 24550 27212 24556
rect 27710 24576 27712 24585
rect 27764 24576 27766 24585
rect 27172 24138 27200 24550
rect 27710 24511 27766 24520
rect 27160 24132 27212 24138
rect 27160 24074 27212 24080
rect 27712 24064 27764 24070
rect 27712 24006 27764 24012
rect 27724 23905 27752 24006
rect 27710 23896 27766 23905
rect 27710 23831 27766 23840
rect 27528 23724 27580 23730
rect 27528 23666 27580 23672
rect 27540 23322 27568 23666
rect 27712 23520 27764 23526
rect 27712 23462 27764 23468
rect 27528 23316 27580 23322
rect 27528 23258 27580 23264
rect 27724 23225 27752 23462
rect 27710 23216 27766 23225
rect 27710 23151 27766 23160
rect 27710 22536 27766 22545
rect 27710 22471 27712 22480
rect 27764 22471 27766 22480
rect 27712 22442 27764 22448
rect 26976 21888 27028 21894
rect 26976 21830 27028 21836
rect 27160 21548 27212 21554
rect 27160 21490 27212 21496
rect 26976 21412 27028 21418
rect 26804 21372 26976 21400
rect 26976 21354 27028 21360
rect 26608 20868 26660 20874
rect 26608 20810 26660 20816
rect 26240 20596 26292 20602
rect 26240 20538 26292 20544
rect 26252 20466 26280 20538
rect 26148 20460 26200 20466
rect 26148 20402 26200 20408
rect 26240 20460 26292 20466
rect 26240 20402 26292 20408
rect 25964 19916 26016 19922
rect 25964 19858 26016 19864
rect 25976 19802 26004 19858
rect 25872 19780 25924 19786
rect 25976 19774 26096 19802
rect 26620 19786 26648 20810
rect 26988 20534 27016 21354
rect 26976 20528 27028 20534
rect 26976 20470 27028 20476
rect 27172 20058 27200 21490
rect 27160 20052 27212 20058
rect 27160 19994 27212 20000
rect 25872 19722 25924 19728
rect 26068 18766 26096 19774
rect 26608 19780 26660 19786
rect 26608 19722 26660 19728
rect 26056 18760 26108 18766
rect 26108 18708 26188 18714
rect 26056 18702 26188 18708
rect 26068 18686 26188 18702
rect 26620 18698 26648 19722
rect 27620 19508 27672 19514
rect 27620 19450 27672 19456
rect 27632 19145 27660 19450
rect 27804 19372 27856 19378
rect 27804 19314 27856 19320
rect 27618 19136 27674 19145
rect 27618 19071 27674 19080
rect 27816 18970 27844 19314
rect 27804 18964 27856 18970
rect 27804 18906 27856 18912
rect 25596 18624 25648 18630
rect 25596 18566 25648 18572
rect 25502 17232 25558 17241
rect 25502 17167 25558 17176
rect 25516 16794 25544 17167
rect 25504 16788 25556 16794
rect 25504 16730 25556 16736
rect 25516 16182 25544 16730
rect 25608 16574 25636 18566
rect 26160 17746 26188 18686
rect 26608 18692 26660 18698
rect 26608 18634 26660 18640
rect 26148 17740 26200 17746
rect 26148 17682 26200 17688
rect 26160 16658 26188 17682
rect 26148 16652 26200 16658
rect 26148 16594 26200 16600
rect 25608 16546 25728 16574
rect 25700 16250 25728 16546
rect 26608 16516 26660 16522
rect 26608 16458 26660 16464
rect 25688 16244 25740 16250
rect 25688 16186 25740 16192
rect 25504 16176 25556 16182
rect 25504 16118 25556 16124
rect 25412 14612 25464 14618
rect 25412 14554 25464 14560
rect 25136 14476 25188 14482
rect 25136 14418 25188 14424
rect 24952 14272 25004 14278
rect 24952 14214 25004 14220
rect 24964 13462 24992 14214
rect 25228 14000 25280 14006
rect 25056 13960 25228 13988
rect 24952 13456 25004 13462
rect 24952 13398 25004 13404
rect 24860 12980 24912 12986
rect 24860 12922 24912 12928
rect 24308 12640 24360 12646
rect 24308 12582 24360 12588
rect 24136 12406 24256 12434
rect 24044 11762 24164 11778
rect 24044 11756 24176 11762
rect 24044 11750 24124 11756
rect 24124 11698 24176 11704
rect 24032 11552 24084 11558
rect 24032 11494 24084 11500
rect 23940 11280 23992 11286
rect 23940 11222 23992 11228
rect 23940 11144 23992 11150
rect 23940 11086 23992 11092
rect 23848 10804 23900 10810
rect 23848 10746 23900 10752
rect 23756 10736 23808 10742
rect 23952 10690 23980 11086
rect 24044 11014 24072 11494
rect 24032 11008 24084 11014
rect 24032 10950 24084 10956
rect 23756 10678 23808 10684
rect 23860 10662 23980 10690
rect 24044 10674 24072 10950
rect 24136 10742 24164 11698
rect 24228 11642 24256 12406
rect 24320 11762 24348 12582
rect 24676 12096 24728 12102
rect 24676 12038 24728 12044
rect 24400 11824 24452 11830
rect 24400 11766 24452 11772
rect 24308 11756 24360 11762
rect 24308 11698 24360 11704
rect 24228 11614 24348 11642
rect 24216 11076 24268 11082
rect 24216 11018 24268 11024
rect 24124 10736 24176 10742
rect 24124 10678 24176 10684
rect 24032 10668 24084 10674
rect 23664 10532 23716 10538
rect 23664 10474 23716 10480
rect 23860 10470 23888 10662
rect 24032 10610 24084 10616
rect 23848 10464 23900 10470
rect 23848 10406 23900 10412
rect 23572 9988 23624 9994
rect 23572 9930 23624 9936
rect 23388 9172 23440 9178
rect 23388 9114 23440 9120
rect 23388 9036 23440 9042
rect 23388 8978 23440 8984
rect 23400 8566 23428 8978
rect 23388 8560 23440 8566
rect 23388 8502 23440 8508
rect 23296 8492 23348 8498
rect 23296 8434 23348 8440
rect 23308 8378 23336 8434
rect 22940 8362 23336 8378
rect 22928 8356 23336 8362
rect 22980 8350 23336 8356
rect 22928 8298 22980 8304
rect 23400 8022 23428 8502
rect 23584 8498 23612 9930
rect 23664 9376 23716 9382
rect 23664 9318 23716 9324
rect 23676 8974 23704 9318
rect 23664 8968 23716 8974
rect 23664 8910 23716 8916
rect 23756 8900 23808 8906
rect 23756 8842 23808 8848
rect 23572 8492 23624 8498
rect 23572 8434 23624 8440
rect 23480 8356 23532 8362
rect 23480 8298 23532 8304
rect 23388 8016 23440 8022
rect 23388 7958 23440 7964
rect 23492 7954 23520 8298
rect 23480 7948 23532 7954
rect 23480 7890 23532 7896
rect 23296 7812 23348 7818
rect 23296 7754 23348 7760
rect 22744 7744 22796 7750
rect 22742 7712 22744 7721
rect 22796 7712 22798 7721
rect 22742 7647 22798 7656
rect 23308 7546 23336 7754
rect 23296 7540 23348 7546
rect 23296 7482 23348 7488
rect 22468 7404 22520 7410
rect 22468 7346 22520 7352
rect 23388 7404 23440 7410
rect 23388 7346 23440 7352
rect 23480 7404 23532 7410
rect 23584 7392 23612 8434
rect 23768 8090 23796 8842
rect 23756 8084 23808 8090
rect 23756 8026 23808 8032
rect 23768 7886 23796 8026
rect 23860 8022 23888 10406
rect 24032 10056 24084 10062
rect 24032 9998 24084 10004
rect 24044 9586 24072 9998
rect 24032 9580 24084 9586
rect 24032 9522 24084 9528
rect 24032 8968 24084 8974
rect 24032 8910 24084 8916
rect 23940 8832 23992 8838
rect 23940 8774 23992 8780
rect 23952 8566 23980 8774
rect 23940 8560 23992 8566
rect 23940 8502 23992 8508
rect 24044 8430 24072 8910
rect 24136 8906 24164 10678
rect 24228 8974 24256 11018
rect 24216 8968 24268 8974
rect 24216 8910 24268 8916
rect 24124 8900 24176 8906
rect 24124 8842 24176 8848
rect 24032 8424 24084 8430
rect 24032 8366 24084 8372
rect 23848 8016 23900 8022
rect 23848 7958 23900 7964
rect 24136 7886 24164 8842
rect 24216 8832 24268 8838
rect 24216 8774 24268 8780
rect 24228 8634 24256 8774
rect 24216 8628 24268 8634
rect 24216 8570 24268 8576
rect 24320 8294 24348 11614
rect 24412 10742 24440 11766
rect 24492 11688 24544 11694
rect 24492 11630 24544 11636
rect 24504 11354 24532 11630
rect 24492 11348 24544 11354
rect 24492 11290 24544 11296
rect 24688 11218 24716 12038
rect 24860 11756 24912 11762
rect 24860 11698 24912 11704
rect 24872 11354 24900 11698
rect 24860 11348 24912 11354
rect 24860 11290 24912 11296
rect 24676 11212 24728 11218
rect 24676 11154 24728 11160
rect 24492 10804 24544 10810
rect 24492 10746 24544 10752
rect 24400 10736 24452 10742
rect 24400 10678 24452 10684
rect 24412 10470 24440 10678
rect 24400 10464 24452 10470
rect 24400 10406 24452 10412
rect 24504 10266 24532 10746
rect 24584 10668 24636 10674
rect 24584 10610 24636 10616
rect 24492 10260 24544 10266
rect 24492 10202 24544 10208
rect 24596 10062 24624 10610
rect 24688 10130 24716 11154
rect 24872 11098 24900 11290
rect 24780 11082 24900 11098
rect 24768 11076 24900 11082
rect 24820 11070 24900 11076
rect 24768 11018 24820 11024
rect 24768 10532 24820 10538
rect 24768 10474 24820 10480
rect 24780 10266 24808 10474
rect 24768 10260 24820 10266
rect 24768 10202 24820 10208
rect 24676 10124 24728 10130
rect 24676 10066 24728 10072
rect 24584 10056 24636 10062
rect 24584 9998 24636 10004
rect 24596 9586 24624 9998
rect 24584 9580 24636 9586
rect 24584 9522 24636 9528
rect 24872 9466 24900 11070
rect 24952 10464 25004 10470
rect 24952 10406 25004 10412
rect 24964 10198 24992 10406
rect 24952 10192 25004 10198
rect 24952 10134 25004 10140
rect 25056 9994 25084 13960
rect 25228 13942 25280 13948
rect 25136 11892 25188 11898
rect 25136 11834 25188 11840
rect 25148 11082 25176 11834
rect 26620 11762 26648 16458
rect 27804 14408 27856 14414
rect 27802 14376 27804 14385
rect 27856 14376 27858 14385
rect 27802 14311 27858 14320
rect 25688 11756 25740 11762
rect 25688 11698 25740 11704
rect 26608 11756 26660 11762
rect 26608 11698 26660 11704
rect 25136 11076 25188 11082
rect 25136 11018 25188 11024
rect 25044 9988 25096 9994
rect 25044 9930 25096 9936
rect 25056 9722 25084 9930
rect 25136 9920 25188 9926
rect 25136 9862 25188 9868
rect 25044 9716 25096 9722
rect 25044 9658 25096 9664
rect 24872 9438 24992 9466
rect 24860 9376 24912 9382
rect 24860 9318 24912 9324
rect 24768 9036 24820 9042
rect 24768 8978 24820 8984
rect 24308 8288 24360 8294
rect 24308 8230 24360 8236
rect 24320 8022 24348 8230
rect 24308 8016 24360 8022
rect 24308 7958 24360 7964
rect 23756 7880 23808 7886
rect 23756 7822 23808 7828
rect 24124 7880 24176 7886
rect 24124 7822 24176 7828
rect 23756 7744 23808 7750
rect 23756 7686 23808 7692
rect 23768 7478 23796 7686
rect 23756 7472 23808 7478
rect 23756 7414 23808 7420
rect 23532 7364 23612 7392
rect 23480 7346 23532 7352
rect 22376 7268 22428 7274
rect 22376 7210 22428 7216
rect 22480 7002 22508 7346
rect 21548 6996 21600 7002
rect 21548 6938 21600 6944
rect 22468 6996 22520 7002
rect 22468 6938 22520 6944
rect 23400 6798 23428 7346
rect 24320 6798 24348 7958
rect 24780 7954 24808 8978
rect 24872 8974 24900 9318
rect 24860 8968 24912 8974
rect 24860 8910 24912 8916
rect 24872 8634 24900 8910
rect 24964 8838 24992 9438
rect 24952 8832 25004 8838
rect 24952 8774 25004 8780
rect 24860 8628 24912 8634
rect 24860 8570 24912 8576
rect 25056 8498 25084 9658
rect 25148 9178 25176 9862
rect 25136 9172 25188 9178
rect 25136 9114 25188 9120
rect 25044 8492 25096 8498
rect 25044 8434 25096 8440
rect 25056 8090 25084 8434
rect 25044 8084 25096 8090
rect 25044 8026 25096 8032
rect 24768 7948 24820 7954
rect 24768 7890 24820 7896
rect 24780 7546 24808 7890
rect 24768 7540 24820 7546
rect 24768 7482 24820 7488
rect 25056 7478 25084 8026
rect 25700 7886 25728 11698
rect 25688 7880 25740 7886
rect 25688 7822 25740 7828
rect 27712 7880 27764 7886
rect 27712 7822 27764 7828
rect 27620 7812 27672 7818
rect 27620 7754 27672 7760
rect 25044 7472 25096 7478
rect 25044 7414 25096 7420
rect 18696 6792 18748 6798
rect 18696 6734 18748 6740
rect 21456 6792 21508 6798
rect 21456 6734 21508 6740
rect 23388 6792 23440 6798
rect 23388 6734 23440 6740
rect 24308 6792 24360 6798
rect 24308 6734 24360 6740
rect 18604 6452 18656 6458
rect 18604 6394 18656 6400
rect 18708 6390 18736 6734
rect 27632 6458 27660 7754
rect 27620 6452 27672 6458
rect 27620 6394 27672 6400
rect 17040 6384 17092 6390
rect 17040 6326 17092 6332
rect 18696 6384 18748 6390
rect 18696 6326 18748 6332
rect 16488 6316 16540 6322
rect 16488 6258 16540 6264
rect 27724 5914 27752 7822
rect 27804 6316 27856 6322
rect 27804 6258 27856 6264
rect 27816 6225 27844 6258
rect 27802 6216 27858 6225
rect 27802 6151 27858 6160
rect 13268 5908 13320 5914
rect 13268 5850 13320 5856
rect 15476 5908 15528 5914
rect 15476 5850 15528 5856
rect 27712 5908 27764 5914
rect 27712 5850 27764 5856
rect 27804 5704 27856 5710
rect 27804 5646 27856 5652
rect 27816 5545 27844 5646
rect 27802 5536 27858 5545
rect 27802 5471 27858 5480
rect 9048 2746 9352 2774
rect 9324 2650 9352 2746
rect 6092 2644 6144 2650
rect 6092 2586 6144 2592
rect 9312 2644 9364 2650
rect 9312 2586 9364 2592
rect 5816 2440 5868 2446
rect 5816 2382 5868 2388
rect 9036 2440 9088 2446
rect 9036 2382 9088 2388
rect 4874 2204 5182 2213
rect 4874 2202 4880 2204
rect 4936 2202 4960 2204
rect 5016 2202 5040 2204
rect 5096 2202 5120 2204
rect 5176 2202 5182 2204
rect 4936 2150 4938 2202
rect 5118 2150 5120 2202
rect 4874 2148 4880 2150
rect 4936 2148 4960 2150
rect 5016 2148 5040 2150
rect 5096 2148 5120 2150
rect 5176 2148 5182 2150
rect 4874 2139 5182 2148
rect 5828 800 5856 2382
rect 9048 800 9076 2382
rect 5814 0 5870 800
rect 9034 0 9090 800
<< via2 >>
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4880 28314 4936 28316
rect 4960 28314 5016 28316
rect 5040 28314 5096 28316
rect 5120 28314 5176 28316
rect 4880 28262 4926 28314
rect 4926 28262 4936 28314
rect 4960 28262 4990 28314
rect 4990 28262 5002 28314
rect 5002 28262 5016 28314
rect 5040 28262 5054 28314
rect 5054 28262 5066 28314
rect 5066 28262 5096 28314
rect 5120 28262 5130 28314
rect 5130 28262 5176 28314
rect 4880 28260 4936 28262
rect 4960 28260 5016 28262
rect 5040 28260 5096 28262
rect 5120 28260 5176 28262
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 846 23976 902 24032
rect 1490 23160 1546 23216
rect 846 22652 848 22672
rect 848 22652 900 22672
rect 900 22652 902 22672
rect 846 22616 902 22652
rect 846 21972 848 21992
rect 848 21972 900 21992
rect 900 21972 902 21992
rect 846 21936 902 21972
rect 1030 21120 1086 21176
rect 1490 20440 1546 20496
rect 846 19896 902 19952
rect 1398 19080 1454 19136
rect 846 16904 902 16960
rect 1398 15000 1454 15056
rect 1398 13640 1454 13696
rect 846 11756 902 11792
rect 846 11736 848 11756
rect 848 11736 900 11756
rect 900 11736 902 11756
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4880 27226 4936 27228
rect 4960 27226 5016 27228
rect 5040 27226 5096 27228
rect 5120 27226 5176 27228
rect 4880 27174 4926 27226
rect 4926 27174 4936 27226
rect 4960 27174 4990 27226
rect 4990 27174 5002 27226
rect 5002 27174 5016 27226
rect 5040 27174 5054 27226
rect 5054 27174 5066 27226
rect 5066 27174 5096 27226
rect 5120 27174 5130 27226
rect 5130 27174 5176 27226
rect 4880 27172 4936 27174
rect 4960 27172 5016 27174
rect 5040 27172 5096 27174
rect 5120 27172 5176 27174
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4880 26138 4936 26140
rect 4960 26138 5016 26140
rect 5040 26138 5096 26140
rect 5120 26138 5176 26140
rect 4880 26086 4926 26138
rect 4926 26086 4936 26138
rect 4960 26086 4990 26138
rect 4990 26086 5002 26138
rect 5002 26086 5016 26138
rect 5040 26086 5054 26138
rect 5054 26086 5066 26138
rect 5066 26086 5096 26138
rect 5120 26086 5130 26138
rect 5130 26086 5176 26138
rect 4880 26084 4936 26086
rect 4960 26084 5016 26086
rect 5040 26084 5096 26086
rect 5120 26084 5176 26086
rect 10322 26968 10378 27024
rect 4880 25050 4936 25052
rect 4960 25050 5016 25052
rect 5040 25050 5096 25052
rect 5120 25050 5176 25052
rect 4880 24998 4926 25050
rect 4926 24998 4936 25050
rect 4960 24998 4990 25050
rect 4990 24998 5002 25050
rect 5002 24998 5016 25050
rect 5040 24998 5054 25050
rect 5054 24998 5066 25050
rect 5066 24998 5096 25050
rect 5120 24998 5130 25050
rect 5130 24998 5176 25050
rect 4880 24996 4936 24998
rect 4960 24996 5016 24998
rect 5040 24996 5096 24998
rect 5120 24996 5176 24998
rect 4880 23962 4936 23964
rect 4960 23962 5016 23964
rect 5040 23962 5096 23964
rect 5120 23962 5176 23964
rect 4880 23910 4926 23962
rect 4926 23910 4936 23962
rect 4960 23910 4990 23962
rect 4990 23910 5002 23962
rect 5002 23910 5016 23962
rect 5040 23910 5054 23962
rect 5054 23910 5066 23962
rect 5066 23910 5096 23962
rect 5120 23910 5130 23962
rect 5130 23910 5176 23962
rect 4880 23908 4936 23910
rect 4960 23908 5016 23910
rect 5040 23908 5096 23910
rect 5120 23908 5176 23910
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4880 22874 4936 22876
rect 4960 22874 5016 22876
rect 5040 22874 5096 22876
rect 5120 22874 5176 22876
rect 4880 22822 4926 22874
rect 4926 22822 4936 22874
rect 4960 22822 4990 22874
rect 4990 22822 5002 22874
rect 5002 22822 5016 22874
rect 5040 22822 5054 22874
rect 5054 22822 5066 22874
rect 5066 22822 5096 22874
rect 5120 22822 5130 22874
rect 5130 22822 5176 22874
rect 4880 22820 4936 22822
rect 4960 22820 5016 22822
rect 5040 22820 5096 22822
rect 5120 22820 5176 22822
rect 4880 21786 4936 21788
rect 4960 21786 5016 21788
rect 5040 21786 5096 21788
rect 5120 21786 5176 21788
rect 4880 21734 4926 21786
rect 4926 21734 4936 21786
rect 4960 21734 4990 21786
rect 4990 21734 5002 21786
rect 5002 21734 5016 21786
rect 5040 21734 5054 21786
rect 5054 21734 5066 21786
rect 5066 21734 5096 21786
rect 5120 21734 5130 21786
rect 5130 21734 5176 21786
rect 4880 21732 4936 21734
rect 4960 21732 5016 21734
rect 5040 21732 5096 21734
rect 5120 21732 5176 21734
rect 4880 20698 4936 20700
rect 4960 20698 5016 20700
rect 5040 20698 5096 20700
rect 5120 20698 5176 20700
rect 4880 20646 4926 20698
rect 4926 20646 4936 20698
rect 4960 20646 4990 20698
rect 4990 20646 5002 20698
rect 5002 20646 5016 20698
rect 5040 20646 5054 20698
rect 5054 20646 5066 20698
rect 5066 20646 5096 20698
rect 5120 20646 5130 20698
rect 5130 20646 5176 20698
rect 4880 20644 4936 20646
rect 4960 20644 5016 20646
rect 5040 20644 5096 20646
rect 5120 20644 5176 20646
rect 4880 19610 4936 19612
rect 4960 19610 5016 19612
rect 5040 19610 5096 19612
rect 5120 19610 5176 19612
rect 4880 19558 4926 19610
rect 4926 19558 4936 19610
rect 4960 19558 4990 19610
rect 4990 19558 5002 19610
rect 5002 19558 5016 19610
rect 5040 19558 5054 19610
rect 5054 19558 5066 19610
rect 5066 19558 5096 19610
rect 5120 19558 5130 19610
rect 5130 19558 5176 19610
rect 4880 19556 4936 19558
rect 4960 19556 5016 19558
rect 5040 19556 5096 19558
rect 5120 19556 5176 19558
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4880 18522 4936 18524
rect 4960 18522 5016 18524
rect 5040 18522 5096 18524
rect 5120 18522 5176 18524
rect 4880 18470 4926 18522
rect 4926 18470 4936 18522
rect 4960 18470 4990 18522
rect 4990 18470 5002 18522
rect 5002 18470 5016 18522
rect 5040 18470 5054 18522
rect 5054 18470 5066 18522
rect 5066 18470 5096 18522
rect 5120 18470 5130 18522
rect 5130 18470 5176 18522
rect 4880 18468 4936 18470
rect 4960 18468 5016 18470
rect 5040 18468 5096 18470
rect 5120 18468 5176 18470
rect 11058 26988 11114 27024
rect 11058 26968 11060 26988
rect 11060 26968 11112 26988
rect 11112 26968 11114 26988
rect 19982 27004 19984 27024
rect 19984 27004 20036 27024
rect 20036 27004 20038 27024
rect 19982 26968 20038 27004
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4880 17434 4936 17436
rect 4960 17434 5016 17436
rect 5040 17434 5096 17436
rect 5120 17434 5176 17436
rect 4880 17382 4926 17434
rect 4926 17382 4936 17434
rect 4960 17382 4990 17434
rect 4990 17382 5002 17434
rect 5002 17382 5016 17434
rect 5040 17382 5054 17434
rect 5054 17382 5066 17434
rect 5066 17382 5096 17434
rect 5120 17382 5130 17434
rect 5130 17382 5176 17434
rect 4880 17380 4936 17382
rect 4960 17380 5016 17382
rect 5040 17380 5096 17382
rect 5120 17380 5176 17382
rect 4880 16346 4936 16348
rect 4960 16346 5016 16348
rect 5040 16346 5096 16348
rect 5120 16346 5176 16348
rect 4880 16294 4926 16346
rect 4926 16294 4936 16346
rect 4960 16294 4990 16346
rect 4990 16294 5002 16346
rect 5002 16294 5016 16346
rect 5040 16294 5054 16346
rect 5054 16294 5066 16346
rect 5066 16294 5096 16346
rect 5120 16294 5130 16346
rect 5130 16294 5176 16346
rect 4880 16292 4936 16294
rect 4960 16292 5016 16294
rect 5040 16292 5096 16294
rect 5120 16292 5176 16294
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4880 15258 4936 15260
rect 4960 15258 5016 15260
rect 5040 15258 5096 15260
rect 5120 15258 5176 15260
rect 4880 15206 4926 15258
rect 4926 15206 4936 15258
rect 4960 15206 4990 15258
rect 4990 15206 5002 15258
rect 5002 15206 5016 15258
rect 5040 15206 5054 15258
rect 5054 15206 5066 15258
rect 5066 15206 5096 15258
rect 5120 15206 5130 15258
rect 5130 15206 5176 15258
rect 4880 15204 4936 15206
rect 4960 15204 5016 15206
rect 5040 15204 5096 15206
rect 5120 15204 5176 15206
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4880 14170 4936 14172
rect 4960 14170 5016 14172
rect 5040 14170 5096 14172
rect 5120 14170 5176 14172
rect 4880 14118 4926 14170
rect 4926 14118 4936 14170
rect 4960 14118 4990 14170
rect 4990 14118 5002 14170
rect 5002 14118 5016 14170
rect 5040 14118 5054 14170
rect 5054 14118 5066 14170
rect 5066 14118 5096 14170
rect 5120 14118 5130 14170
rect 5130 14118 5176 14170
rect 4880 14116 4936 14118
rect 4960 14116 5016 14118
rect 5040 14116 5096 14118
rect 5120 14116 5176 14118
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4880 13082 4936 13084
rect 4960 13082 5016 13084
rect 5040 13082 5096 13084
rect 5120 13082 5176 13084
rect 4880 13030 4926 13082
rect 4926 13030 4936 13082
rect 4960 13030 4990 13082
rect 4990 13030 5002 13082
rect 5002 13030 5016 13082
rect 5040 13030 5054 13082
rect 5054 13030 5066 13082
rect 5066 13030 5096 13082
rect 5120 13030 5130 13082
rect 5130 13030 5176 13082
rect 4880 13028 4936 13030
rect 4960 13028 5016 13030
rect 5040 13028 5096 13030
rect 5120 13028 5176 13030
rect 4880 11994 4936 11996
rect 4960 11994 5016 11996
rect 5040 11994 5096 11996
rect 5120 11994 5176 11996
rect 4880 11942 4926 11994
rect 4926 11942 4936 11994
rect 4960 11942 4990 11994
rect 4990 11942 5002 11994
rect 5002 11942 5016 11994
rect 5040 11942 5054 11994
rect 5054 11942 5066 11994
rect 5066 11942 5096 11994
rect 5120 11942 5130 11994
rect 5130 11942 5176 11994
rect 4880 11940 4936 11942
rect 4960 11940 5016 11942
rect 5040 11940 5096 11942
rect 5120 11940 5176 11942
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4880 10906 4936 10908
rect 4960 10906 5016 10908
rect 5040 10906 5096 10908
rect 5120 10906 5176 10908
rect 4880 10854 4926 10906
rect 4926 10854 4936 10906
rect 4960 10854 4990 10906
rect 4990 10854 5002 10906
rect 5002 10854 5016 10906
rect 5040 10854 5054 10906
rect 5054 10854 5066 10906
rect 5066 10854 5096 10906
rect 5120 10854 5130 10906
rect 5130 10854 5176 10906
rect 4880 10852 4936 10854
rect 4960 10852 5016 10854
rect 5040 10852 5096 10854
rect 5120 10852 5176 10854
rect 4880 9818 4936 9820
rect 4960 9818 5016 9820
rect 5040 9818 5096 9820
rect 5120 9818 5176 9820
rect 4880 9766 4926 9818
rect 4926 9766 4936 9818
rect 4960 9766 4990 9818
rect 4990 9766 5002 9818
rect 5002 9766 5016 9818
rect 5040 9766 5054 9818
rect 5054 9766 5066 9818
rect 5066 9766 5096 9818
rect 5120 9766 5130 9818
rect 5130 9766 5176 9818
rect 4880 9764 4936 9766
rect 4960 9764 5016 9766
rect 5040 9764 5096 9766
rect 5120 9764 5176 9766
rect 4880 8730 4936 8732
rect 4960 8730 5016 8732
rect 5040 8730 5096 8732
rect 5120 8730 5176 8732
rect 4880 8678 4926 8730
rect 4926 8678 4936 8730
rect 4960 8678 4990 8730
rect 4990 8678 5002 8730
rect 5002 8678 5016 8730
rect 5040 8678 5054 8730
rect 5054 8678 5066 8730
rect 5066 8678 5096 8730
rect 5120 8678 5130 8730
rect 5130 8678 5176 8730
rect 4880 8676 4936 8678
rect 4960 8676 5016 8678
rect 5040 8676 5096 8678
rect 5120 8676 5176 8678
rect 4880 7642 4936 7644
rect 4960 7642 5016 7644
rect 5040 7642 5096 7644
rect 5120 7642 5176 7644
rect 4880 7590 4926 7642
rect 4926 7590 4936 7642
rect 4960 7590 4990 7642
rect 4990 7590 5002 7642
rect 5002 7590 5016 7642
rect 5040 7590 5054 7642
rect 5054 7590 5066 7642
rect 5066 7590 5096 7642
rect 5120 7590 5130 7642
rect 5130 7590 5176 7642
rect 4880 7588 4936 7590
rect 4960 7588 5016 7590
rect 5040 7588 5096 7590
rect 5120 7588 5176 7590
rect 11794 20848 11850 20904
rect 20626 26988 20682 27024
rect 20626 26968 20628 26988
rect 20628 26968 20680 26988
rect 20680 26968 20682 26988
rect 22282 27004 22284 27024
rect 22284 27004 22336 27024
rect 22336 27004 22338 27024
rect 22282 26968 22338 27004
rect 12530 20748 12532 20768
rect 12532 20748 12584 20768
rect 12584 20748 12586 20768
rect 12530 20712 12586 20748
rect 12530 20476 12532 20496
rect 12532 20476 12584 20496
rect 12584 20476 12586 20496
rect 12530 20440 12586 20476
rect 12898 21548 12954 21584
rect 12898 21528 12900 21548
rect 12900 21528 12952 21548
rect 12952 21528 12954 21548
rect 10046 12960 10102 13016
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4880 6554 4936 6556
rect 4960 6554 5016 6556
rect 5040 6554 5096 6556
rect 5120 6554 5176 6556
rect 4880 6502 4926 6554
rect 4926 6502 4936 6554
rect 4960 6502 4990 6554
rect 4990 6502 5002 6554
rect 5002 6502 5016 6554
rect 5040 6502 5054 6554
rect 5054 6502 5066 6554
rect 5066 6502 5096 6554
rect 5120 6502 5130 6554
rect 5130 6502 5176 6554
rect 4880 6500 4936 6502
rect 4960 6500 5016 6502
rect 5040 6500 5096 6502
rect 5120 6500 5176 6502
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4880 5466 4936 5468
rect 4960 5466 5016 5468
rect 5040 5466 5096 5468
rect 5120 5466 5176 5468
rect 4880 5414 4926 5466
rect 4926 5414 4936 5466
rect 4960 5414 4990 5466
rect 4990 5414 5002 5466
rect 5002 5414 5016 5466
rect 5040 5414 5054 5466
rect 5054 5414 5066 5466
rect 5066 5414 5096 5466
rect 5120 5414 5130 5466
rect 5130 5414 5176 5466
rect 4880 5412 4936 5414
rect 4960 5412 5016 5414
rect 5040 5412 5096 5414
rect 5120 5412 5176 5414
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4880 4378 4936 4380
rect 4960 4378 5016 4380
rect 5040 4378 5096 4380
rect 5120 4378 5176 4380
rect 4880 4326 4926 4378
rect 4926 4326 4936 4378
rect 4960 4326 4990 4378
rect 4990 4326 5002 4378
rect 5002 4326 5016 4378
rect 5040 4326 5054 4378
rect 5054 4326 5066 4378
rect 5066 4326 5096 4378
rect 5120 4326 5130 4378
rect 5130 4326 5176 4378
rect 4880 4324 4936 4326
rect 4960 4324 5016 4326
rect 5040 4324 5096 4326
rect 5120 4324 5176 4326
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4880 3290 4936 3292
rect 4960 3290 5016 3292
rect 5040 3290 5096 3292
rect 5120 3290 5176 3292
rect 4880 3238 4926 3290
rect 4926 3238 4936 3290
rect 4960 3238 4990 3290
rect 4990 3238 5002 3290
rect 5002 3238 5016 3290
rect 5040 3238 5054 3290
rect 5054 3238 5066 3290
rect 5066 3238 5096 3290
rect 5120 3238 5130 3290
rect 5130 3238 5176 3290
rect 4880 3236 4936 3238
rect 4960 3236 5016 3238
rect 5040 3236 5096 3238
rect 5120 3236 5176 3238
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 11334 11620 11390 11656
rect 11334 11600 11336 11620
rect 11336 11600 11388 11620
rect 11388 11600 11390 11620
rect 13634 21548 13690 21584
rect 13634 21528 13636 21548
rect 13636 21528 13688 21548
rect 13688 21528 13690 21548
rect 13450 20032 13506 20088
rect 13910 20304 13966 20360
rect 14186 20884 14188 20904
rect 14188 20884 14240 20904
rect 14240 20884 14242 20904
rect 14186 20848 14242 20884
rect 14094 20476 14096 20496
rect 14096 20476 14148 20496
rect 14148 20476 14150 20496
rect 14094 20440 14150 20476
rect 11702 13912 11758 13968
rect 13542 14456 13598 14512
rect 11978 11092 11980 11112
rect 11980 11092 12032 11112
rect 12032 11092 12034 11112
rect 11978 11056 12034 11092
rect 13542 13640 13598 13696
rect 12990 11892 13046 11928
rect 12990 11872 12992 11892
rect 12992 11872 13044 11892
rect 13044 11872 13046 11892
rect 12898 11056 12954 11112
rect 12162 7792 12218 7848
rect 12714 9444 12770 9480
rect 12714 9424 12716 9444
rect 12716 9424 12768 9444
rect 12768 9424 12770 9444
rect 12162 7540 12218 7576
rect 12162 7520 12164 7540
rect 12164 7520 12216 7540
rect 12216 7520 12218 7540
rect 12622 7112 12678 7168
rect 16946 24132 17002 24168
rect 16946 24112 16948 24132
rect 16948 24112 17000 24132
rect 17000 24112 17002 24132
rect 13174 8084 13230 8120
rect 13174 8064 13176 8084
rect 13176 8064 13228 8084
rect 13228 8064 13230 8084
rect 12898 6740 12900 6760
rect 12900 6740 12952 6760
rect 12952 6740 12954 6760
rect 12898 6704 12954 6740
rect 14186 7656 14242 7712
rect 13266 6976 13322 7032
rect 13910 7248 13966 7304
rect 14830 7404 14886 7440
rect 14830 7384 14832 7404
rect 14832 7384 14884 7404
rect 14884 7384 14886 7404
rect 14278 7248 14334 7304
rect 15842 19352 15898 19408
rect 15842 17196 15898 17232
rect 15842 17176 15844 17196
rect 15844 17176 15896 17196
rect 15896 17176 15898 17196
rect 17314 21528 17370 21584
rect 15934 17040 15990 17096
rect 15566 11892 15622 11928
rect 15566 11872 15568 11892
rect 15568 11872 15620 11892
rect 15620 11872 15622 11892
rect 15934 13776 15990 13832
rect 15842 12960 15898 13016
rect 16210 17040 16266 17096
rect 16670 16632 16726 16688
rect 17314 20324 17370 20360
rect 17314 20304 17316 20324
rect 17316 20304 17368 20324
rect 17368 20304 17370 20324
rect 16946 17620 16948 17640
rect 16948 17620 17000 17640
rect 17000 17620 17002 17640
rect 16946 17584 17002 17620
rect 15566 11056 15622 11112
rect 15934 11056 15990 11112
rect 15474 10648 15530 10704
rect 15290 8064 15346 8120
rect 15382 7404 15438 7440
rect 15382 7384 15384 7404
rect 15384 7384 15436 7404
rect 15436 7384 15438 7404
rect 15014 6996 15070 7032
rect 15014 6976 15016 6996
rect 15016 6976 15068 6996
rect 15068 6976 15070 6996
rect 16302 11056 16358 11112
rect 15842 7792 15898 7848
rect 15934 7112 15990 7168
rect 16210 7792 16266 7848
rect 16118 6976 16174 7032
rect 16762 11872 16818 11928
rect 17222 17040 17278 17096
rect 18050 24112 18106 24168
rect 18050 16532 18052 16552
rect 18052 16532 18104 16552
rect 18104 16532 18106 16552
rect 18050 16496 18106 16532
rect 17038 12008 17094 12064
rect 18050 13912 18106 13968
rect 17498 10668 17554 10704
rect 17498 10648 17500 10668
rect 17500 10648 17552 10668
rect 17552 10648 17554 10668
rect 16946 10004 16948 10024
rect 16948 10004 17000 10024
rect 17000 10004 17002 10024
rect 16946 9968 17002 10004
rect 16578 7520 16634 7576
rect 16578 7248 16634 7304
rect 17958 9968 18014 10024
rect 17222 8200 17278 8256
rect 17130 7928 17186 7984
rect 17774 7828 17776 7848
rect 17776 7828 17828 7848
rect 17828 7828 17830 7848
rect 17774 7792 17830 7828
rect 19154 20324 19210 20360
rect 19154 20304 19156 20324
rect 19156 20304 19208 20324
rect 19208 20304 19210 20324
rect 19062 17584 19118 17640
rect 19062 17040 19118 17096
rect 18326 10004 18328 10024
rect 18328 10004 18380 10024
rect 18380 10004 18382 10024
rect 18326 9968 18382 10004
rect 18602 7828 18604 7848
rect 18604 7828 18656 7848
rect 18656 7828 18658 7848
rect 17498 7112 17554 7168
rect 18602 7792 18658 7828
rect 18878 7928 18934 7984
rect 18786 7384 18842 7440
rect 19798 21292 19800 21312
rect 19800 21292 19852 21312
rect 19852 21292 19854 21312
rect 19798 21256 19854 21292
rect 24582 26968 24638 27024
rect 24950 26988 25006 27024
rect 24950 26968 24952 26988
rect 24952 26968 25004 26988
rect 25004 26968 25006 26988
rect 25318 27532 25374 27568
rect 25318 27512 25320 27532
rect 25320 27512 25372 27532
rect 25372 27512 25374 27532
rect 20534 17332 20590 17368
rect 20534 17312 20536 17332
rect 20536 17312 20588 17332
rect 20588 17312 20590 17332
rect 22742 20304 22798 20360
rect 19522 13776 19578 13832
rect 19706 12844 19762 12880
rect 19706 12824 19708 12844
rect 19708 12824 19760 12844
rect 19760 12824 19762 12844
rect 20810 17196 20866 17232
rect 20810 17176 20812 17196
rect 20812 17176 20864 17196
rect 20864 17176 20866 17196
rect 21270 16632 21326 16688
rect 21822 17312 21878 17368
rect 22466 19372 22522 19408
rect 22466 19352 22468 19372
rect 22468 19352 22520 19372
rect 22520 19352 22522 19372
rect 20534 15272 20590 15328
rect 20626 13812 20628 13832
rect 20628 13812 20680 13832
rect 20680 13812 20682 13832
rect 20074 11600 20130 11656
rect 20626 13776 20682 13812
rect 20902 13776 20958 13832
rect 19614 8200 19670 8256
rect 19522 7828 19524 7848
rect 19524 7828 19576 7848
rect 19576 7828 19578 7848
rect 19522 7792 19578 7828
rect 20074 8084 20130 8120
rect 20074 8064 20076 8084
rect 20076 8064 20128 8084
rect 20128 8064 20130 8084
rect 20074 7540 20130 7576
rect 20074 7520 20076 7540
rect 20076 7520 20128 7540
rect 20128 7520 20130 7540
rect 20994 7928 21050 7984
rect 20902 7404 20958 7440
rect 20902 7384 20904 7404
rect 20904 7384 20956 7404
rect 20956 7384 20958 7404
rect 22282 14456 22338 14512
rect 22282 13776 22338 13832
rect 21822 12824 21878 12880
rect 23938 21256 23994 21312
rect 25134 22888 25190 22944
rect 25870 26988 25926 27024
rect 25870 26968 25872 26988
rect 25872 26968 25924 26988
rect 25924 26968 25926 26988
rect 26330 27532 26386 27568
rect 26330 27512 26332 27532
rect 26332 27512 26384 27532
rect 26384 27512 26386 27532
rect 22558 9580 22614 9616
rect 22558 9560 22560 9580
rect 22560 9560 22612 9580
rect 22612 9560 22614 9580
rect 22374 9460 22376 9480
rect 22376 9460 22428 9480
rect 22428 9460 22430 9480
rect 22374 9424 22430 9460
rect 22282 7792 22338 7848
rect 22190 7520 22246 7576
rect 24030 15444 24032 15464
rect 24032 15444 24084 15464
rect 24084 15444 24086 15464
rect 24030 15408 24086 15444
rect 24582 13268 24584 13288
rect 24584 13268 24636 13288
rect 24636 13268 24638 13288
rect 24582 13232 24638 13268
rect 27710 25880 27766 25936
rect 27710 25200 27766 25256
rect 27710 24556 27712 24576
rect 27712 24556 27764 24576
rect 27764 24556 27766 24576
rect 27710 24520 27766 24556
rect 27710 23840 27766 23896
rect 27710 23160 27766 23216
rect 27710 22500 27766 22536
rect 27710 22480 27712 22500
rect 27712 22480 27764 22500
rect 27764 22480 27766 22500
rect 27618 19080 27674 19136
rect 25502 17176 25558 17232
rect 22742 7692 22744 7712
rect 22744 7692 22796 7712
rect 22796 7692 22798 7712
rect 22742 7656 22798 7692
rect 27802 14356 27804 14376
rect 27804 14356 27856 14376
rect 27856 14356 27858 14376
rect 27802 14320 27858 14356
rect 27802 6160 27858 6216
rect 27802 5480 27858 5536
rect 4880 2202 4936 2204
rect 4960 2202 5016 2204
rect 5040 2202 5096 2204
rect 5120 2202 5176 2204
rect 4880 2150 4926 2202
rect 4926 2150 4936 2202
rect 4960 2150 4990 2202
rect 4990 2150 5002 2202
rect 5002 2150 5016 2202
rect 5040 2150 5054 2202
rect 5054 2150 5066 2202
rect 5066 2150 5096 2202
rect 5120 2150 5130 2202
rect 5130 2150 5176 2202
rect 4880 2148 4936 2150
rect 4960 2148 5016 2150
rect 5040 2148 5096 2150
rect 5120 2148 5176 2150
<< metal3 >>
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 4870 28320 5186 28321
rect 4870 28256 4876 28320
rect 4940 28256 4956 28320
rect 5020 28256 5036 28320
rect 5100 28256 5116 28320
rect 5180 28256 5186 28320
rect 4870 28255 5186 28256
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 25313 27570 25379 27573
rect 26325 27570 26391 27573
rect 25313 27568 26391 27570
rect 25313 27512 25318 27568
rect 25374 27512 26330 27568
rect 26386 27512 26391 27568
rect 25313 27510 26391 27512
rect 25313 27507 25379 27510
rect 26325 27507 26391 27510
rect 4870 27232 5186 27233
rect 4870 27168 4876 27232
rect 4940 27168 4956 27232
rect 5020 27168 5036 27232
rect 5100 27168 5116 27232
rect 5180 27168 5186 27232
rect 4870 27167 5186 27168
rect 10317 27026 10383 27029
rect 11053 27026 11119 27029
rect 10317 27024 11119 27026
rect 10317 26968 10322 27024
rect 10378 26968 11058 27024
rect 11114 26968 11119 27024
rect 10317 26966 11119 26968
rect 10317 26963 10383 26966
rect 11053 26963 11119 26966
rect 19977 27026 20043 27029
rect 20621 27026 20687 27029
rect 19977 27024 20687 27026
rect 19977 26968 19982 27024
rect 20038 26968 20626 27024
rect 20682 26968 20687 27024
rect 19977 26966 20687 26968
rect 19977 26963 20043 26966
rect 20621 26963 20687 26966
rect 22277 27026 22343 27029
rect 24577 27026 24643 27029
rect 22277 27024 24643 27026
rect 22277 26968 22282 27024
rect 22338 26968 24582 27024
rect 24638 26968 24643 27024
rect 22277 26966 24643 26968
rect 22277 26963 22343 26966
rect 24577 26963 24643 26966
rect 24945 27026 25011 27029
rect 25865 27026 25931 27029
rect 24945 27024 25931 27026
rect 24945 26968 24950 27024
rect 25006 26968 25870 27024
rect 25926 26968 25931 27024
rect 24945 26966 25931 26968
rect 24945 26963 25011 26966
rect 25865 26963 25931 26966
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 4870 26144 5186 26145
rect 4870 26080 4876 26144
rect 4940 26080 4956 26144
rect 5020 26080 5036 26144
rect 5100 26080 5116 26144
rect 5180 26080 5186 26144
rect 4870 26079 5186 26080
rect 27705 25938 27771 25941
rect 28532 25938 29332 25968
rect 27705 25936 29332 25938
rect 27705 25880 27710 25936
rect 27766 25880 29332 25936
rect 27705 25878 29332 25880
rect 27705 25875 27771 25878
rect 28532 25848 29332 25878
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 27705 25258 27771 25261
rect 28532 25258 29332 25288
rect 27705 25256 29332 25258
rect 27705 25200 27710 25256
rect 27766 25200 29332 25256
rect 27705 25198 29332 25200
rect 27705 25195 27771 25198
rect 28532 25168 29332 25198
rect 4870 25056 5186 25057
rect 4870 24992 4876 25056
rect 4940 24992 4956 25056
rect 5020 24992 5036 25056
rect 5100 24992 5116 25056
rect 5180 24992 5186 25056
rect 4870 24991 5186 24992
rect 27705 24578 27771 24581
rect 28532 24578 29332 24608
rect 27705 24576 29332 24578
rect 27705 24520 27710 24576
rect 27766 24520 29332 24576
rect 27705 24518 29332 24520
rect 27705 24515 27771 24518
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 28532 24488 29332 24518
rect 4210 24447 4526 24448
rect 16941 24170 17007 24173
rect 18045 24170 18111 24173
rect 16941 24168 18111 24170
rect 16941 24112 16946 24168
rect 17002 24112 18050 24168
rect 18106 24112 18111 24168
rect 16941 24110 18111 24112
rect 16941 24107 17007 24110
rect 18045 24107 18111 24110
rect 841 24034 907 24037
rect 798 24032 907 24034
rect 798 23976 846 24032
rect 902 23976 907 24032
rect 798 23971 907 23976
rect 798 23928 858 23971
rect 0 23838 858 23928
rect 4870 23968 5186 23969
rect 4870 23904 4876 23968
rect 4940 23904 4956 23968
rect 5020 23904 5036 23968
rect 5100 23904 5116 23968
rect 5180 23904 5186 23968
rect 4870 23903 5186 23904
rect 27705 23898 27771 23901
rect 28532 23898 29332 23928
rect 27705 23896 29332 23898
rect 27705 23840 27710 23896
rect 27766 23840 29332 23896
rect 27705 23838 29332 23840
rect 0 23808 800 23838
rect 27705 23835 27771 23838
rect 28532 23808 29332 23838
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 0 23218 800 23248
rect 1485 23218 1551 23221
rect 0 23216 1551 23218
rect 0 23160 1490 23216
rect 1546 23160 1551 23216
rect 0 23158 1551 23160
rect 0 23128 800 23158
rect 1485 23155 1551 23158
rect 27705 23218 27771 23221
rect 28532 23218 29332 23248
rect 27705 23216 29332 23218
rect 27705 23160 27710 23216
rect 27766 23160 29332 23216
rect 27705 23158 29332 23160
rect 27705 23155 27771 23158
rect 28532 23128 29332 23158
rect 24894 22884 24900 22948
rect 24964 22946 24970 22948
rect 25129 22946 25195 22949
rect 24964 22944 25195 22946
rect 24964 22888 25134 22944
rect 25190 22888 25195 22944
rect 24964 22886 25195 22888
rect 24964 22884 24970 22886
rect 25129 22883 25195 22886
rect 4870 22880 5186 22881
rect 4870 22816 4876 22880
rect 4940 22816 4956 22880
rect 5020 22816 5036 22880
rect 5100 22816 5116 22880
rect 5180 22816 5186 22880
rect 4870 22815 5186 22816
rect 841 22674 907 22677
rect 798 22672 907 22674
rect 798 22616 846 22672
rect 902 22616 907 22672
rect 798 22611 907 22616
rect 798 22568 858 22611
rect 0 22478 858 22568
rect 27705 22538 27771 22541
rect 28532 22538 29332 22568
rect 27705 22536 29332 22538
rect 27705 22480 27710 22536
rect 27766 22480 29332 22536
rect 27705 22478 29332 22480
rect 0 22448 800 22478
rect 27705 22475 27771 22478
rect 28532 22448 29332 22478
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 841 21994 907 21997
rect 798 21992 907 21994
rect 798 21936 846 21992
rect 902 21936 907 21992
rect 798 21931 907 21936
rect 798 21888 858 21931
rect 0 21798 858 21888
rect 0 21768 800 21798
rect 4870 21792 5186 21793
rect 4870 21728 4876 21792
rect 4940 21728 4956 21792
rect 5020 21728 5036 21792
rect 5100 21728 5116 21792
rect 5180 21728 5186 21792
rect 4870 21727 5186 21728
rect 12893 21586 12959 21589
rect 13629 21586 13695 21589
rect 17309 21586 17375 21589
rect 12893 21584 17375 21586
rect 12893 21528 12898 21584
rect 12954 21528 13634 21584
rect 13690 21528 17314 21584
rect 17370 21528 17375 21584
rect 12893 21526 17375 21528
rect 12893 21523 12959 21526
rect 13629 21523 13695 21526
rect 17309 21523 17375 21526
rect 19793 21314 19859 21317
rect 23933 21314 23999 21317
rect 19793 21312 23999 21314
rect 19793 21256 19798 21312
rect 19854 21256 23938 21312
rect 23994 21256 23999 21312
rect 19793 21254 23999 21256
rect 19793 21251 19859 21254
rect 23933 21251 23999 21254
rect 4210 21248 4526 21249
rect 0 21178 800 21208
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 1025 21178 1091 21181
rect 0 21176 1091 21178
rect 0 21120 1030 21176
rect 1086 21120 1091 21176
rect 0 21118 1091 21120
rect 0 21088 800 21118
rect 1025 21115 1091 21118
rect 11789 20906 11855 20909
rect 14181 20906 14247 20909
rect 11789 20904 14247 20906
rect 11789 20848 11794 20904
rect 11850 20848 14186 20904
rect 14242 20848 14247 20904
rect 11789 20846 14247 20848
rect 11789 20843 11855 20846
rect 14181 20843 14247 20846
rect 12525 20772 12591 20773
rect 12525 20770 12572 20772
rect 12480 20768 12572 20770
rect 12480 20712 12530 20768
rect 12480 20710 12572 20712
rect 12525 20708 12572 20710
rect 12636 20708 12642 20772
rect 12525 20707 12591 20708
rect 4870 20704 5186 20705
rect 4870 20640 4876 20704
rect 4940 20640 4956 20704
rect 5020 20640 5036 20704
rect 5100 20640 5116 20704
rect 5180 20640 5186 20704
rect 4870 20639 5186 20640
rect 0 20498 800 20528
rect 1485 20498 1551 20501
rect 0 20496 1551 20498
rect 0 20440 1490 20496
rect 1546 20440 1551 20496
rect 0 20438 1551 20440
rect 0 20408 800 20438
rect 1485 20435 1551 20438
rect 12525 20498 12591 20501
rect 14089 20498 14155 20501
rect 12525 20496 14155 20498
rect 12525 20440 12530 20496
rect 12586 20440 14094 20496
rect 14150 20440 14155 20496
rect 12525 20438 14155 20440
rect 12525 20435 12591 20438
rect 14089 20435 14155 20438
rect 13905 20362 13971 20365
rect 17309 20362 17375 20365
rect 19149 20362 19215 20365
rect 22737 20362 22803 20365
rect 13905 20360 17375 20362
rect 13905 20304 13910 20360
rect 13966 20304 17314 20360
rect 17370 20304 17375 20360
rect 13905 20302 17375 20304
rect 13905 20299 13971 20302
rect 17309 20299 17375 20302
rect 17910 20360 22803 20362
rect 17910 20304 19154 20360
rect 19210 20304 22742 20360
rect 22798 20304 22803 20360
rect 17910 20302 22803 20304
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 13445 20090 13511 20093
rect 17910 20090 17970 20302
rect 19149 20299 19215 20302
rect 22737 20299 22803 20302
rect 13445 20088 17970 20090
rect 13445 20032 13450 20088
rect 13506 20032 17970 20088
rect 13445 20030 17970 20032
rect 13445 20027 13511 20030
rect 841 19954 907 19957
rect 798 19952 907 19954
rect 798 19896 846 19952
rect 902 19896 907 19952
rect 798 19891 907 19896
rect 798 19848 858 19891
rect 0 19758 858 19848
rect 0 19728 800 19758
rect 4870 19616 5186 19617
rect 4870 19552 4876 19616
rect 4940 19552 4956 19616
rect 5020 19552 5036 19616
rect 5100 19552 5116 19616
rect 5180 19552 5186 19616
rect 4870 19551 5186 19552
rect 15837 19410 15903 19413
rect 22461 19410 22527 19413
rect 15837 19408 22527 19410
rect 15837 19352 15842 19408
rect 15898 19352 22466 19408
rect 22522 19352 22527 19408
rect 15837 19350 22527 19352
rect 15837 19347 15903 19350
rect 22461 19347 22527 19350
rect 0 19138 800 19168
rect 1393 19138 1459 19141
rect 0 19136 1459 19138
rect 0 19080 1398 19136
rect 1454 19080 1459 19136
rect 0 19078 1459 19080
rect 0 19048 800 19078
rect 1393 19075 1459 19078
rect 27613 19138 27679 19141
rect 28532 19138 29332 19168
rect 27613 19136 29332 19138
rect 27613 19080 27618 19136
rect 27674 19080 29332 19136
rect 27613 19078 29332 19080
rect 27613 19075 27679 19078
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 28532 19048 29332 19078
rect 4210 19007 4526 19008
rect 4870 18528 5186 18529
rect 4870 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5186 18528
rect 4870 18463 5186 18464
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 16941 17642 17007 17645
rect 19057 17642 19123 17645
rect 16941 17640 19123 17642
rect 16941 17584 16946 17640
rect 17002 17584 19062 17640
rect 19118 17584 19123 17640
rect 16941 17582 19123 17584
rect 16941 17579 17007 17582
rect 19057 17579 19123 17582
rect 4870 17440 5186 17441
rect 4870 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5186 17440
rect 4870 17375 5186 17376
rect 20529 17370 20595 17373
rect 21817 17370 21883 17373
rect 20529 17368 21883 17370
rect 20529 17312 20534 17368
rect 20590 17312 21822 17368
rect 21878 17312 21883 17368
rect 20529 17310 21883 17312
rect 20529 17307 20595 17310
rect 21817 17307 21883 17310
rect 15837 17234 15903 17237
rect 20805 17234 20871 17237
rect 24894 17234 24900 17236
rect 15837 17232 20871 17234
rect 15837 17176 15842 17232
rect 15898 17176 20810 17232
rect 20866 17176 20871 17232
rect 15837 17174 20871 17176
rect 15837 17171 15903 17174
rect 20805 17171 20871 17174
rect 22050 17174 24900 17234
rect 0 17098 800 17128
rect 15929 17098 15995 17101
rect 16205 17098 16271 17101
rect 17217 17098 17283 17101
rect 0 17008 858 17098
rect 15929 17096 17283 17098
rect 15929 17040 15934 17096
rect 15990 17040 16210 17096
rect 16266 17040 17222 17096
rect 17278 17040 17283 17096
rect 15929 17038 17283 17040
rect 15929 17035 15995 17038
rect 16205 17035 16271 17038
rect 17217 17035 17283 17038
rect 19057 17098 19123 17101
rect 22050 17098 22110 17174
rect 24894 17172 24900 17174
rect 24964 17234 24970 17236
rect 25497 17234 25563 17237
rect 24964 17232 25563 17234
rect 24964 17176 25502 17232
rect 25558 17176 25563 17232
rect 24964 17174 25563 17176
rect 24964 17172 24970 17174
rect 25497 17171 25563 17174
rect 19057 17096 22110 17098
rect 19057 17040 19062 17096
rect 19118 17040 22110 17096
rect 19057 17038 22110 17040
rect 19057 17035 19123 17038
rect 798 16965 858 17008
rect 798 16960 907 16965
rect 798 16904 846 16960
rect 902 16904 907 16960
rect 798 16902 907 16904
rect 841 16899 907 16902
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 16665 16690 16731 16693
rect 21265 16690 21331 16693
rect 16665 16688 21331 16690
rect 16665 16632 16670 16688
rect 16726 16632 21270 16688
rect 21326 16632 21331 16688
rect 16665 16630 21331 16632
rect 16665 16627 16731 16630
rect 21265 16627 21331 16630
rect 18045 16554 18111 16557
rect 19190 16554 19196 16556
rect 18045 16552 19196 16554
rect 18045 16496 18050 16552
rect 18106 16496 19196 16552
rect 18045 16494 19196 16496
rect 18045 16491 18111 16494
rect 19190 16492 19196 16494
rect 19260 16492 19266 16556
rect 4870 16352 5186 16353
rect 4870 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5186 16352
rect 4870 16287 5186 16288
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 24025 15468 24091 15469
rect 23974 15404 23980 15468
rect 24044 15466 24091 15468
rect 24044 15464 24136 15466
rect 24086 15408 24136 15464
rect 24044 15406 24136 15408
rect 24044 15404 24091 15406
rect 24025 15403 24091 15404
rect 20529 15332 20595 15333
rect 20478 15330 20484 15332
rect 20438 15270 20484 15330
rect 20548 15328 20595 15332
rect 20590 15272 20595 15328
rect 20478 15268 20484 15270
rect 20548 15268 20595 15272
rect 20529 15267 20595 15268
rect 4870 15264 5186 15265
rect 4870 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5186 15264
rect 4870 15199 5186 15200
rect 0 15058 800 15088
rect 1393 15058 1459 15061
rect 0 15056 1459 15058
rect 0 15000 1398 15056
rect 1454 15000 1459 15056
rect 0 14998 1459 15000
rect 0 14968 800 14998
rect 1393 14995 1459 14998
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 13537 14514 13603 14517
rect 22277 14514 22343 14517
rect 13537 14512 22343 14514
rect 13537 14456 13542 14512
rect 13598 14456 22282 14512
rect 22338 14456 22343 14512
rect 13537 14454 22343 14456
rect 13537 14451 13603 14454
rect 22277 14451 22343 14454
rect 27797 14378 27863 14381
rect 28532 14378 29332 14408
rect 27797 14376 29332 14378
rect 27797 14320 27802 14376
rect 27858 14320 29332 14376
rect 27797 14318 29332 14320
rect 27797 14315 27863 14318
rect 28532 14288 29332 14318
rect 4870 14176 5186 14177
rect 4870 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5186 14176
rect 4870 14111 5186 14112
rect 11697 13970 11763 13973
rect 18045 13970 18111 13973
rect 11697 13968 18111 13970
rect 11697 13912 11702 13968
rect 11758 13912 18050 13968
rect 18106 13912 18111 13968
rect 11697 13910 18111 13912
rect 11697 13907 11763 13910
rect 18045 13907 18111 13910
rect 15929 13834 15995 13837
rect 19517 13834 19583 13837
rect 20621 13834 20687 13837
rect 15929 13832 20687 13834
rect 15929 13776 15934 13832
rect 15990 13776 19522 13832
rect 19578 13776 20626 13832
rect 20682 13776 20687 13832
rect 15929 13774 20687 13776
rect 15929 13771 15995 13774
rect 19517 13771 19583 13774
rect 20621 13771 20687 13774
rect 20897 13834 20963 13837
rect 22277 13834 22343 13837
rect 20897 13832 22343 13834
rect 20897 13776 20902 13832
rect 20958 13776 22282 13832
rect 22338 13776 22343 13832
rect 20897 13774 22343 13776
rect 20897 13771 20963 13774
rect 22277 13771 22343 13774
rect 0 13698 800 13728
rect 1393 13698 1459 13701
rect 0 13696 1459 13698
rect 0 13640 1398 13696
rect 1454 13640 1459 13696
rect 0 13638 1459 13640
rect 0 13608 800 13638
rect 1393 13635 1459 13638
rect 12566 13636 12572 13700
rect 12636 13698 12642 13700
rect 13537 13698 13603 13701
rect 12636 13696 13603 13698
rect 12636 13640 13542 13696
rect 13598 13640 13603 13696
rect 12636 13638 13603 13640
rect 12636 13636 12642 13638
rect 13537 13635 13603 13638
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 24577 13292 24643 13293
rect 24526 13228 24532 13292
rect 24596 13290 24643 13292
rect 24596 13288 24688 13290
rect 24638 13232 24688 13288
rect 24596 13230 24688 13232
rect 24596 13228 24643 13230
rect 24577 13227 24643 13228
rect 4870 13088 5186 13089
rect 4870 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5186 13088
rect 4870 13023 5186 13024
rect 10041 13018 10107 13021
rect 15837 13018 15903 13021
rect 10041 13016 15903 13018
rect 10041 12960 10046 13016
rect 10102 12960 15842 13016
rect 15898 12960 15903 13016
rect 10041 12958 15903 12960
rect 10041 12955 10107 12958
rect 15837 12955 15903 12958
rect 19701 12882 19767 12885
rect 21817 12882 21883 12885
rect 19701 12880 21883 12882
rect 19701 12824 19706 12880
rect 19762 12824 21822 12880
rect 21878 12824 21883 12880
rect 19701 12822 21883 12824
rect 19701 12819 19767 12822
rect 21817 12819 21883 12822
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 17033 12066 17099 12069
rect 12988 12064 17099 12066
rect 12988 12008 17038 12064
rect 17094 12008 17099 12064
rect 12988 12006 17099 12008
rect 4870 12000 5186 12001
rect 4870 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5186 12000
rect 4870 11935 5186 11936
rect 12988 11933 13048 12006
rect 17033 12003 17099 12006
rect 12750 11868 12756 11932
rect 12820 11930 12826 11932
rect 12985 11930 13051 11933
rect 12820 11928 13051 11930
rect 12820 11872 12990 11928
rect 13046 11872 13051 11928
rect 12820 11870 13051 11872
rect 12820 11868 12826 11870
rect 12985 11867 13051 11870
rect 15561 11930 15627 11933
rect 16757 11930 16823 11933
rect 15561 11928 16823 11930
rect 15561 11872 15566 11928
rect 15622 11872 16762 11928
rect 16818 11872 16823 11928
rect 15561 11870 16823 11872
rect 15561 11867 15627 11870
rect 16757 11867 16823 11870
rect 841 11794 907 11797
rect 798 11792 907 11794
rect 798 11736 846 11792
rect 902 11736 907 11792
rect 798 11731 907 11736
rect 798 11688 858 11731
rect 0 11598 858 11688
rect 11329 11658 11395 11661
rect 20069 11658 20135 11661
rect 11329 11656 20135 11658
rect 11329 11600 11334 11656
rect 11390 11600 20074 11656
rect 20130 11600 20135 11656
rect 11329 11598 20135 11600
rect 0 11568 800 11598
rect 11329 11595 11395 11598
rect 20069 11595 20135 11598
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 11973 11114 12039 11117
rect 12893 11114 12959 11117
rect 11973 11112 12959 11114
rect 11973 11056 11978 11112
rect 12034 11056 12898 11112
rect 12954 11056 12959 11112
rect 11973 11054 12959 11056
rect 11973 11051 12039 11054
rect 12893 11051 12959 11054
rect 15561 11114 15627 11117
rect 15929 11114 15995 11117
rect 16297 11114 16363 11117
rect 15561 11112 16363 11114
rect 15561 11056 15566 11112
rect 15622 11056 15934 11112
rect 15990 11056 16302 11112
rect 16358 11056 16363 11112
rect 15561 11054 16363 11056
rect 15561 11051 15627 11054
rect 15929 11051 15995 11054
rect 16297 11051 16363 11054
rect 4870 10912 5186 10913
rect 4870 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5186 10912
rect 4870 10847 5186 10848
rect 15469 10706 15535 10709
rect 17493 10706 17559 10709
rect 15469 10704 17559 10706
rect 15469 10648 15474 10704
rect 15530 10648 17498 10704
rect 17554 10648 17559 10704
rect 15469 10646 17559 10648
rect 15469 10643 15535 10646
rect 17493 10643 17559 10646
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 16941 10026 17007 10029
rect 17953 10026 18019 10029
rect 18321 10026 18387 10029
rect 16941 10024 18387 10026
rect 16941 9968 16946 10024
rect 17002 9968 17958 10024
rect 18014 9968 18326 10024
rect 18382 9968 18387 10024
rect 16941 9966 18387 9968
rect 16941 9963 17007 9966
rect 17953 9963 18019 9966
rect 18321 9963 18387 9966
rect 4870 9824 5186 9825
rect 4870 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5186 9824
rect 4870 9759 5186 9760
rect 22553 9618 22619 9621
rect 24526 9618 24532 9620
rect 22553 9616 24532 9618
rect 22553 9560 22558 9616
rect 22614 9560 24532 9616
rect 22553 9558 24532 9560
rect 22553 9555 22619 9558
rect 24526 9556 24532 9558
rect 24596 9556 24602 9620
rect 12709 9484 12775 9485
rect 12709 9482 12756 9484
rect 12664 9480 12756 9482
rect 12664 9424 12714 9480
rect 12664 9422 12756 9424
rect 12709 9420 12756 9422
rect 12820 9420 12826 9484
rect 22369 9482 22435 9485
rect 23974 9482 23980 9484
rect 22369 9480 23980 9482
rect 22369 9424 22374 9480
rect 22430 9424 23980 9480
rect 22369 9422 23980 9424
rect 12709 9419 12775 9420
rect 22369 9419 22435 9422
rect 23974 9420 23980 9422
rect 24044 9420 24050 9484
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 4870 8736 5186 8737
rect 4870 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5186 8736
rect 4870 8671 5186 8672
rect 17217 8258 17283 8261
rect 19609 8258 19675 8261
rect 17217 8256 19675 8258
rect 17217 8200 17222 8256
rect 17278 8200 19614 8256
rect 19670 8200 19675 8256
rect 17217 8198 19675 8200
rect 17217 8195 17283 8198
rect 19609 8195 19675 8198
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 13169 8122 13235 8125
rect 15285 8122 15351 8125
rect 13169 8120 15351 8122
rect 13169 8064 13174 8120
rect 13230 8064 15290 8120
rect 15346 8064 15351 8120
rect 13169 8062 15351 8064
rect 13169 8059 13235 8062
rect 15285 8059 15351 8062
rect 19190 8060 19196 8124
rect 19260 8122 19266 8124
rect 20069 8122 20135 8125
rect 19260 8120 20135 8122
rect 19260 8064 20074 8120
rect 20130 8064 20135 8120
rect 19260 8062 20135 8064
rect 19260 8060 19266 8062
rect 20069 8059 20135 8062
rect 17125 7986 17191 7989
rect 18873 7986 18939 7989
rect 20989 7986 21055 7989
rect 16070 7984 21055 7986
rect 16070 7928 17130 7984
rect 17186 7928 18878 7984
rect 18934 7928 20994 7984
rect 21050 7928 21055 7984
rect 16070 7926 21055 7928
rect 12157 7850 12223 7853
rect 15837 7850 15903 7853
rect 16070 7850 16130 7926
rect 17125 7923 17191 7926
rect 18873 7923 18939 7926
rect 20989 7923 21055 7926
rect 12157 7848 16130 7850
rect 12157 7792 12162 7848
rect 12218 7792 15842 7848
rect 15898 7792 16130 7848
rect 12157 7790 16130 7792
rect 16205 7850 16271 7853
rect 17769 7850 17835 7853
rect 18597 7850 18663 7853
rect 16205 7848 18663 7850
rect 16205 7792 16210 7848
rect 16266 7792 17774 7848
rect 17830 7792 18602 7848
rect 18658 7792 18663 7848
rect 16205 7790 18663 7792
rect 12157 7787 12223 7790
rect 15837 7787 15903 7790
rect 16205 7787 16271 7790
rect 17769 7787 17835 7790
rect 18597 7787 18663 7790
rect 19517 7850 19583 7853
rect 22277 7850 22343 7853
rect 19517 7848 22343 7850
rect 19517 7792 19522 7848
rect 19578 7792 22282 7848
rect 22338 7792 22343 7848
rect 19517 7790 22343 7792
rect 19517 7787 19583 7790
rect 22277 7787 22343 7790
rect 14181 7714 14247 7717
rect 22737 7714 22803 7717
rect 14181 7712 22803 7714
rect 14181 7656 14186 7712
rect 14242 7656 22742 7712
rect 22798 7656 22803 7712
rect 14181 7654 22803 7656
rect 14181 7651 14247 7654
rect 22737 7651 22803 7654
rect 4870 7648 5186 7649
rect 4870 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5186 7648
rect 4870 7583 5186 7584
rect 12157 7578 12223 7581
rect 16573 7578 16639 7581
rect 12157 7576 16639 7578
rect 12157 7520 12162 7576
rect 12218 7520 16578 7576
rect 16634 7520 16639 7576
rect 12157 7518 16639 7520
rect 12157 7515 12223 7518
rect 16573 7515 16639 7518
rect 20069 7578 20135 7581
rect 22185 7578 22251 7581
rect 20069 7576 22251 7578
rect 20069 7520 20074 7576
rect 20130 7520 22190 7576
rect 22246 7520 22251 7576
rect 20069 7518 22251 7520
rect 20069 7515 20135 7518
rect 22185 7515 22251 7518
rect 14825 7442 14891 7445
rect 15377 7442 15443 7445
rect 14825 7440 15443 7442
rect 14825 7384 14830 7440
rect 14886 7384 15382 7440
rect 15438 7384 15443 7440
rect 14825 7382 15443 7384
rect 14825 7379 14891 7382
rect 15377 7379 15443 7382
rect 18781 7442 18847 7445
rect 20897 7442 20963 7445
rect 18781 7440 20963 7442
rect 18781 7384 18786 7440
rect 18842 7384 20902 7440
rect 20958 7384 20963 7440
rect 18781 7382 20963 7384
rect 18781 7379 18847 7382
rect 20897 7379 20963 7382
rect 13905 7306 13971 7309
rect 14273 7306 14339 7309
rect 16573 7306 16639 7309
rect 13905 7304 16639 7306
rect 13905 7248 13910 7304
rect 13966 7248 14278 7304
rect 14334 7248 16578 7304
rect 16634 7248 16639 7304
rect 13905 7246 16639 7248
rect 13905 7243 13971 7246
rect 14273 7243 14339 7246
rect 16573 7243 16639 7246
rect 12617 7170 12683 7173
rect 15929 7170 15995 7173
rect 17493 7170 17559 7173
rect 12617 7168 17559 7170
rect 12617 7112 12622 7168
rect 12678 7112 15934 7168
rect 15990 7112 17498 7168
rect 17554 7112 17559 7168
rect 12617 7110 17559 7112
rect 12617 7107 12683 7110
rect 15929 7107 15995 7110
rect 17493 7107 17559 7110
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 13261 7034 13327 7037
rect 15009 7034 15075 7037
rect 16113 7034 16179 7037
rect 13261 7032 16179 7034
rect 13261 6976 13266 7032
rect 13322 6976 15014 7032
rect 15070 6976 16118 7032
rect 16174 6976 16179 7032
rect 13261 6974 16179 6976
rect 13261 6971 13327 6974
rect 15009 6971 15075 6974
rect 16113 6971 16179 6974
rect 12750 6700 12756 6764
rect 12820 6762 12826 6764
rect 12893 6762 12959 6765
rect 12820 6760 12959 6762
rect 12820 6704 12898 6760
rect 12954 6704 12959 6760
rect 12820 6702 12959 6704
rect 12820 6700 12826 6702
rect 12893 6699 12959 6702
rect 4870 6560 5186 6561
rect 4870 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5186 6560
rect 4870 6495 5186 6496
rect 27797 6218 27863 6221
rect 28532 6218 29332 6248
rect 27797 6216 29332 6218
rect 27797 6160 27802 6216
rect 27858 6160 29332 6216
rect 27797 6158 29332 6160
rect 27797 6155 27863 6158
rect 28532 6128 29332 6158
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 27797 5538 27863 5541
rect 28532 5538 29332 5568
rect 27797 5536 29332 5538
rect 27797 5480 27802 5536
rect 27858 5480 29332 5536
rect 27797 5478 29332 5480
rect 27797 5475 27863 5478
rect 4870 5472 5186 5473
rect 4870 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5186 5472
rect 28532 5448 29332 5478
rect 4870 5407 5186 5408
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 20478 4796 20484 4860
rect 20548 4858 20554 4860
rect 28532 4858 29332 4888
rect 20548 4798 29332 4858
rect 20548 4796 20554 4798
rect 28532 4768 29332 4798
rect 4870 4384 5186 4385
rect 4870 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5186 4384
rect 4870 4319 5186 4320
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 4870 3296 5186 3297
rect 4870 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5186 3296
rect 4870 3231 5186 3232
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 4870 2208 5186 2209
rect 4870 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5186 2208
rect 4870 2143 5186 2144
<< via3 >>
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 4876 28316 4940 28320
rect 4876 28260 4880 28316
rect 4880 28260 4936 28316
rect 4936 28260 4940 28316
rect 4876 28256 4940 28260
rect 4956 28316 5020 28320
rect 4956 28260 4960 28316
rect 4960 28260 5016 28316
rect 5016 28260 5020 28316
rect 4956 28256 5020 28260
rect 5036 28316 5100 28320
rect 5036 28260 5040 28316
rect 5040 28260 5096 28316
rect 5096 28260 5100 28316
rect 5036 28256 5100 28260
rect 5116 28316 5180 28320
rect 5116 28260 5120 28316
rect 5120 28260 5176 28316
rect 5176 28260 5180 28316
rect 5116 28256 5180 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 4876 27228 4940 27232
rect 4876 27172 4880 27228
rect 4880 27172 4936 27228
rect 4936 27172 4940 27228
rect 4876 27168 4940 27172
rect 4956 27228 5020 27232
rect 4956 27172 4960 27228
rect 4960 27172 5016 27228
rect 5016 27172 5020 27228
rect 4956 27168 5020 27172
rect 5036 27228 5100 27232
rect 5036 27172 5040 27228
rect 5040 27172 5096 27228
rect 5096 27172 5100 27228
rect 5036 27168 5100 27172
rect 5116 27228 5180 27232
rect 5116 27172 5120 27228
rect 5120 27172 5176 27228
rect 5176 27172 5180 27228
rect 5116 27168 5180 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 4876 26140 4940 26144
rect 4876 26084 4880 26140
rect 4880 26084 4936 26140
rect 4936 26084 4940 26140
rect 4876 26080 4940 26084
rect 4956 26140 5020 26144
rect 4956 26084 4960 26140
rect 4960 26084 5016 26140
rect 5016 26084 5020 26140
rect 4956 26080 5020 26084
rect 5036 26140 5100 26144
rect 5036 26084 5040 26140
rect 5040 26084 5096 26140
rect 5096 26084 5100 26140
rect 5036 26080 5100 26084
rect 5116 26140 5180 26144
rect 5116 26084 5120 26140
rect 5120 26084 5176 26140
rect 5176 26084 5180 26140
rect 5116 26080 5180 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 4876 25052 4940 25056
rect 4876 24996 4880 25052
rect 4880 24996 4936 25052
rect 4936 24996 4940 25052
rect 4876 24992 4940 24996
rect 4956 25052 5020 25056
rect 4956 24996 4960 25052
rect 4960 24996 5016 25052
rect 5016 24996 5020 25052
rect 4956 24992 5020 24996
rect 5036 25052 5100 25056
rect 5036 24996 5040 25052
rect 5040 24996 5096 25052
rect 5096 24996 5100 25052
rect 5036 24992 5100 24996
rect 5116 25052 5180 25056
rect 5116 24996 5120 25052
rect 5120 24996 5176 25052
rect 5176 24996 5180 25052
rect 5116 24992 5180 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 4876 23964 4940 23968
rect 4876 23908 4880 23964
rect 4880 23908 4936 23964
rect 4936 23908 4940 23964
rect 4876 23904 4940 23908
rect 4956 23964 5020 23968
rect 4956 23908 4960 23964
rect 4960 23908 5016 23964
rect 5016 23908 5020 23964
rect 4956 23904 5020 23908
rect 5036 23964 5100 23968
rect 5036 23908 5040 23964
rect 5040 23908 5096 23964
rect 5096 23908 5100 23964
rect 5036 23904 5100 23908
rect 5116 23964 5180 23968
rect 5116 23908 5120 23964
rect 5120 23908 5176 23964
rect 5176 23908 5180 23964
rect 5116 23904 5180 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 24900 22884 24964 22948
rect 4876 22876 4940 22880
rect 4876 22820 4880 22876
rect 4880 22820 4936 22876
rect 4936 22820 4940 22876
rect 4876 22816 4940 22820
rect 4956 22876 5020 22880
rect 4956 22820 4960 22876
rect 4960 22820 5016 22876
rect 5016 22820 5020 22876
rect 4956 22816 5020 22820
rect 5036 22876 5100 22880
rect 5036 22820 5040 22876
rect 5040 22820 5096 22876
rect 5096 22820 5100 22876
rect 5036 22816 5100 22820
rect 5116 22876 5180 22880
rect 5116 22820 5120 22876
rect 5120 22820 5176 22876
rect 5176 22820 5180 22876
rect 5116 22816 5180 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 4876 21788 4940 21792
rect 4876 21732 4880 21788
rect 4880 21732 4936 21788
rect 4936 21732 4940 21788
rect 4876 21728 4940 21732
rect 4956 21788 5020 21792
rect 4956 21732 4960 21788
rect 4960 21732 5016 21788
rect 5016 21732 5020 21788
rect 4956 21728 5020 21732
rect 5036 21788 5100 21792
rect 5036 21732 5040 21788
rect 5040 21732 5096 21788
rect 5096 21732 5100 21788
rect 5036 21728 5100 21732
rect 5116 21788 5180 21792
rect 5116 21732 5120 21788
rect 5120 21732 5176 21788
rect 5176 21732 5180 21788
rect 5116 21728 5180 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 12572 20768 12636 20772
rect 12572 20712 12586 20768
rect 12586 20712 12636 20768
rect 12572 20708 12636 20712
rect 4876 20700 4940 20704
rect 4876 20644 4880 20700
rect 4880 20644 4936 20700
rect 4936 20644 4940 20700
rect 4876 20640 4940 20644
rect 4956 20700 5020 20704
rect 4956 20644 4960 20700
rect 4960 20644 5016 20700
rect 5016 20644 5020 20700
rect 4956 20640 5020 20644
rect 5036 20700 5100 20704
rect 5036 20644 5040 20700
rect 5040 20644 5096 20700
rect 5096 20644 5100 20700
rect 5036 20640 5100 20644
rect 5116 20700 5180 20704
rect 5116 20644 5120 20700
rect 5120 20644 5176 20700
rect 5176 20644 5180 20700
rect 5116 20640 5180 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 4876 19612 4940 19616
rect 4876 19556 4880 19612
rect 4880 19556 4936 19612
rect 4936 19556 4940 19612
rect 4876 19552 4940 19556
rect 4956 19612 5020 19616
rect 4956 19556 4960 19612
rect 4960 19556 5016 19612
rect 5016 19556 5020 19612
rect 4956 19552 5020 19556
rect 5036 19612 5100 19616
rect 5036 19556 5040 19612
rect 5040 19556 5096 19612
rect 5096 19556 5100 19612
rect 5036 19552 5100 19556
rect 5116 19612 5180 19616
rect 5116 19556 5120 19612
rect 5120 19556 5176 19612
rect 5176 19556 5180 19612
rect 5116 19552 5180 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 4876 18524 4940 18528
rect 4876 18468 4880 18524
rect 4880 18468 4936 18524
rect 4936 18468 4940 18524
rect 4876 18464 4940 18468
rect 4956 18524 5020 18528
rect 4956 18468 4960 18524
rect 4960 18468 5016 18524
rect 5016 18468 5020 18524
rect 4956 18464 5020 18468
rect 5036 18524 5100 18528
rect 5036 18468 5040 18524
rect 5040 18468 5096 18524
rect 5096 18468 5100 18524
rect 5036 18464 5100 18468
rect 5116 18524 5180 18528
rect 5116 18468 5120 18524
rect 5120 18468 5176 18524
rect 5176 18468 5180 18524
rect 5116 18464 5180 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 4876 17436 4940 17440
rect 4876 17380 4880 17436
rect 4880 17380 4936 17436
rect 4936 17380 4940 17436
rect 4876 17376 4940 17380
rect 4956 17436 5020 17440
rect 4956 17380 4960 17436
rect 4960 17380 5016 17436
rect 5016 17380 5020 17436
rect 4956 17376 5020 17380
rect 5036 17436 5100 17440
rect 5036 17380 5040 17436
rect 5040 17380 5096 17436
rect 5096 17380 5100 17436
rect 5036 17376 5100 17380
rect 5116 17436 5180 17440
rect 5116 17380 5120 17436
rect 5120 17380 5176 17436
rect 5176 17380 5180 17436
rect 5116 17376 5180 17380
rect 24900 17172 24964 17236
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 19196 16492 19260 16556
rect 4876 16348 4940 16352
rect 4876 16292 4880 16348
rect 4880 16292 4936 16348
rect 4936 16292 4940 16348
rect 4876 16288 4940 16292
rect 4956 16348 5020 16352
rect 4956 16292 4960 16348
rect 4960 16292 5016 16348
rect 5016 16292 5020 16348
rect 4956 16288 5020 16292
rect 5036 16348 5100 16352
rect 5036 16292 5040 16348
rect 5040 16292 5096 16348
rect 5096 16292 5100 16348
rect 5036 16288 5100 16292
rect 5116 16348 5180 16352
rect 5116 16292 5120 16348
rect 5120 16292 5176 16348
rect 5176 16292 5180 16348
rect 5116 16288 5180 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 23980 15464 24044 15468
rect 23980 15408 24030 15464
rect 24030 15408 24044 15464
rect 23980 15404 24044 15408
rect 20484 15328 20548 15332
rect 20484 15272 20534 15328
rect 20534 15272 20548 15328
rect 20484 15268 20548 15272
rect 4876 15260 4940 15264
rect 4876 15204 4880 15260
rect 4880 15204 4936 15260
rect 4936 15204 4940 15260
rect 4876 15200 4940 15204
rect 4956 15260 5020 15264
rect 4956 15204 4960 15260
rect 4960 15204 5016 15260
rect 5016 15204 5020 15260
rect 4956 15200 5020 15204
rect 5036 15260 5100 15264
rect 5036 15204 5040 15260
rect 5040 15204 5096 15260
rect 5096 15204 5100 15260
rect 5036 15200 5100 15204
rect 5116 15260 5180 15264
rect 5116 15204 5120 15260
rect 5120 15204 5176 15260
rect 5176 15204 5180 15260
rect 5116 15200 5180 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 4876 14172 4940 14176
rect 4876 14116 4880 14172
rect 4880 14116 4936 14172
rect 4936 14116 4940 14172
rect 4876 14112 4940 14116
rect 4956 14172 5020 14176
rect 4956 14116 4960 14172
rect 4960 14116 5016 14172
rect 5016 14116 5020 14172
rect 4956 14112 5020 14116
rect 5036 14172 5100 14176
rect 5036 14116 5040 14172
rect 5040 14116 5096 14172
rect 5096 14116 5100 14172
rect 5036 14112 5100 14116
rect 5116 14172 5180 14176
rect 5116 14116 5120 14172
rect 5120 14116 5176 14172
rect 5176 14116 5180 14172
rect 5116 14112 5180 14116
rect 12572 13636 12636 13700
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 24532 13288 24596 13292
rect 24532 13232 24582 13288
rect 24582 13232 24596 13288
rect 24532 13228 24596 13232
rect 4876 13084 4940 13088
rect 4876 13028 4880 13084
rect 4880 13028 4936 13084
rect 4936 13028 4940 13084
rect 4876 13024 4940 13028
rect 4956 13084 5020 13088
rect 4956 13028 4960 13084
rect 4960 13028 5016 13084
rect 5016 13028 5020 13084
rect 4956 13024 5020 13028
rect 5036 13084 5100 13088
rect 5036 13028 5040 13084
rect 5040 13028 5096 13084
rect 5096 13028 5100 13084
rect 5036 13024 5100 13028
rect 5116 13084 5180 13088
rect 5116 13028 5120 13084
rect 5120 13028 5176 13084
rect 5176 13028 5180 13084
rect 5116 13024 5180 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 4876 11996 4940 12000
rect 4876 11940 4880 11996
rect 4880 11940 4936 11996
rect 4936 11940 4940 11996
rect 4876 11936 4940 11940
rect 4956 11996 5020 12000
rect 4956 11940 4960 11996
rect 4960 11940 5016 11996
rect 5016 11940 5020 11996
rect 4956 11936 5020 11940
rect 5036 11996 5100 12000
rect 5036 11940 5040 11996
rect 5040 11940 5096 11996
rect 5096 11940 5100 11996
rect 5036 11936 5100 11940
rect 5116 11996 5180 12000
rect 5116 11940 5120 11996
rect 5120 11940 5176 11996
rect 5176 11940 5180 11996
rect 5116 11936 5180 11940
rect 12756 11868 12820 11932
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 4876 10908 4940 10912
rect 4876 10852 4880 10908
rect 4880 10852 4936 10908
rect 4936 10852 4940 10908
rect 4876 10848 4940 10852
rect 4956 10908 5020 10912
rect 4956 10852 4960 10908
rect 4960 10852 5016 10908
rect 5016 10852 5020 10908
rect 4956 10848 5020 10852
rect 5036 10908 5100 10912
rect 5036 10852 5040 10908
rect 5040 10852 5096 10908
rect 5096 10852 5100 10908
rect 5036 10848 5100 10852
rect 5116 10908 5180 10912
rect 5116 10852 5120 10908
rect 5120 10852 5176 10908
rect 5176 10852 5180 10908
rect 5116 10848 5180 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 4876 9820 4940 9824
rect 4876 9764 4880 9820
rect 4880 9764 4936 9820
rect 4936 9764 4940 9820
rect 4876 9760 4940 9764
rect 4956 9820 5020 9824
rect 4956 9764 4960 9820
rect 4960 9764 5016 9820
rect 5016 9764 5020 9820
rect 4956 9760 5020 9764
rect 5036 9820 5100 9824
rect 5036 9764 5040 9820
rect 5040 9764 5096 9820
rect 5096 9764 5100 9820
rect 5036 9760 5100 9764
rect 5116 9820 5180 9824
rect 5116 9764 5120 9820
rect 5120 9764 5176 9820
rect 5176 9764 5180 9820
rect 5116 9760 5180 9764
rect 24532 9556 24596 9620
rect 12756 9480 12820 9484
rect 12756 9424 12770 9480
rect 12770 9424 12820 9480
rect 12756 9420 12820 9424
rect 23980 9420 24044 9484
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 4876 8732 4940 8736
rect 4876 8676 4880 8732
rect 4880 8676 4936 8732
rect 4936 8676 4940 8732
rect 4876 8672 4940 8676
rect 4956 8732 5020 8736
rect 4956 8676 4960 8732
rect 4960 8676 5016 8732
rect 5016 8676 5020 8732
rect 4956 8672 5020 8676
rect 5036 8732 5100 8736
rect 5036 8676 5040 8732
rect 5040 8676 5096 8732
rect 5096 8676 5100 8732
rect 5036 8672 5100 8676
rect 5116 8732 5180 8736
rect 5116 8676 5120 8732
rect 5120 8676 5176 8732
rect 5176 8676 5180 8732
rect 5116 8672 5180 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 19196 8060 19260 8124
rect 4876 7644 4940 7648
rect 4876 7588 4880 7644
rect 4880 7588 4936 7644
rect 4936 7588 4940 7644
rect 4876 7584 4940 7588
rect 4956 7644 5020 7648
rect 4956 7588 4960 7644
rect 4960 7588 5016 7644
rect 5016 7588 5020 7644
rect 4956 7584 5020 7588
rect 5036 7644 5100 7648
rect 5036 7588 5040 7644
rect 5040 7588 5096 7644
rect 5096 7588 5100 7644
rect 5036 7584 5100 7588
rect 5116 7644 5180 7648
rect 5116 7588 5120 7644
rect 5120 7588 5176 7644
rect 5176 7588 5180 7644
rect 5116 7584 5180 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 12756 6700 12820 6764
rect 4876 6556 4940 6560
rect 4876 6500 4880 6556
rect 4880 6500 4936 6556
rect 4936 6500 4940 6556
rect 4876 6496 4940 6500
rect 4956 6556 5020 6560
rect 4956 6500 4960 6556
rect 4960 6500 5016 6556
rect 5016 6500 5020 6556
rect 4956 6496 5020 6500
rect 5036 6556 5100 6560
rect 5036 6500 5040 6556
rect 5040 6500 5096 6556
rect 5096 6500 5100 6556
rect 5036 6496 5100 6500
rect 5116 6556 5180 6560
rect 5116 6500 5120 6556
rect 5120 6500 5176 6556
rect 5176 6500 5180 6556
rect 5116 6496 5180 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 4876 5468 4940 5472
rect 4876 5412 4880 5468
rect 4880 5412 4936 5468
rect 4936 5412 4940 5468
rect 4876 5408 4940 5412
rect 4956 5468 5020 5472
rect 4956 5412 4960 5468
rect 4960 5412 5016 5468
rect 5016 5412 5020 5468
rect 4956 5408 5020 5412
rect 5036 5468 5100 5472
rect 5036 5412 5040 5468
rect 5040 5412 5096 5468
rect 5096 5412 5100 5468
rect 5036 5408 5100 5412
rect 5116 5468 5180 5472
rect 5116 5412 5120 5468
rect 5120 5412 5176 5468
rect 5176 5412 5180 5468
rect 5116 5408 5180 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 20484 4796 20548 4860
rect 4876 4380 4940 4384
rect 4876 4324 4880 4380
rect 4880 4324 4936 4380
rect 4936 4324 4940 4380
rect 4876 4320 4940 4324
rect 4956 4380 5020 4384
rect 4956 4324 4960 4380
rect 4960 4324 5016 4380
rect 5016 4324 5020 4380
rect 4956 4320 5020 4324
rect 5036 4380 5100 4384
rect 5036 4324 5040 4380
rect 5040 4324 5096 4380
rect 5096 4324 5100 4380
rect 5036 4320 5100 4324
rect 5116 4380 5180 4384
rect 5116 4324 5120 4380
rect 5120 4324 5176 4380
rect 5176 4324 5180 4380
rect 5116 4320 5180 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 4876 3292 4940 3296
rect 4876 3236 4880 3292
rect 4880 3236 4936 3292
rect 4936 3236 4940 3292
rect 4876 3232 4940 3236
rect 4956 3292 5020 3296
rect 4956 3236 4960 3292
rect 4960 3236 5016 3292
rect 5016 3236 5020 3292
rect 4956 3232 5020 3236
rect 5036 3292 5100 3296
rect 5036 3236 5040 3292
rect 5040 3236 5096 3292
rect 5096 3236 5100 3292
rect 5036 3232 5100 3236
rect 5116 3292 5180 3296
rect 5116 3236 5120 3292
rect 5120 3236 5176 3292
rect 5176 3236 5180 3292
rect 5116 3232 5180 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 4876 2204 4940 2208
rect 4876 2148 4880 2204
rect 4880 2148 4936 2204
rect 4936 2148 4940 2204
rect 4876 2144 4940 2148
rect 4956 2204 5020 2208
rect 4956 2148 4960 2204
rect 4960 2148 5016 2204
rect 5016 2148 5020 2204
rect 4956 2144 5020 2148
rect 5036 2204 5100 2208
rect 5036 2148 5040 2204
rect 5040 2148 5096 2204
rect 5096 2148 5100 2204
rect 5036 2144 5100 2148
rect 5116 2204 5180 2208
rect 5116 2148 5120 2204
rect 5120 2148 5176 2204
rect 5176 2148 5180 2204
rect 5116 2144 5180 2148
<< metal4 >>
rect 4208 28864 4528 28880
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 4868 28320 5188 28880
rect 4868 28256 4876 28320
rect 4940 28256 4956 28320
rect 5020 28256 5036 28320
rect 5100 28256 5116 28320
rect 5180 28256 5188 28320
rect 4868 27232 5188 28256
rect 4868 27168 4876 27232
rect 4940 27168 4956 27232
rect 5020 27168 5036 27232
rect 5100 27168 5116 27232
rect 5180 27168 5188 27232
rect 4868 26144 5188 27168
rect 4868 26080 4876 26144
rect 4940 26080 4956 26144
rect 5020 26080 5036 26144
rect 5100 26080 5116 26144
rect 5180 26080 5188 26144
rect 4868 25056 5188 26080
rect 4868 24992 4876 25056
rect 4940 24992 4956 25056
rect 5020 24992 5036 25056
rect 5100 24992 5116 25056
rect 5180 24992 5188 25056
rect 4868 23968 5188 24992
rect 4868 23904 4876 23968
rect 4940 23904 4956 23968
rect 5020 23904 5036 23968
rect 5100 23904 5116 23968
rect 5180 23904 5188 23968
rect 4868 22880 5188 23904
rect 24899 22948 24965 22949
rect 24899 22884 24900 22948
rect 24964 22884 24965 22948
rect 24899 22883 24965 22884
rect 4868 22816 4876 22880
rect 4940 22816 4956 22880
rect 5020 22816 5036 22880
rect 5100 22816 5116 22880
rect 5180 22816 5188 22880
rect 4868 21792 5188 22816
rect 4868 21728 4876 21792
rect 4940 21728 4956 21792
rect 5020 21728 5036 21792
rect 5100 21728 5116 21792
rect 5180 21728 5188 21792
rect 4868 20704 5188 21728
rect 12571 20772 12637 20773
rect 12571 20708 12572 20772
rect 12636 20708 12637 20772
rect 12571 20707 12637 20708
rect 4868 20640 4876 20704
rect 4940 20640 4956 20704
rect 5020 20640 5036 20704
rect 5100 20640 5116 20704
rect 5180 20640 5188 20704
rect 4868 19616 5188 20640
rect 4868 19552 4876 19616
rect 4940 19552 4956 19616
rect 5020 19552 5036 19616
rect 5100 19552 5116 19616
rect 5180 19552 5188 19616
rect 4868 18528 5188 19552
rect 4868 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5188 18528
rect 4868 17440 5188 18464
rect 4868 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5188 17440
rect 4868 16352 5188 17376
rect 4868 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5188 16352
rect 4868 15264 5188 16288
rect 4868 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5188 15264
rect 4868 14176 5188 15200
rect 4868 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5188 14176
rect 4868 13088 5188 14112
rect 12574 13701 12634 20707
rect 24902 17237 24962 22883
rect 24899 17236 24965 17237
rect 24899 17172 24900 17236
rect 24964 17172 24965 17236
rect 24899 17171 24965 17172
rect 19195 16556 19261 16557
rect 19195 16492 19196 16556
rect 19260 16492 19261 16556
rect 19195 16491 19261 16492
rect 12571 13700 12637 13701
rect 12571 13636 12572 13700
rect 12636 13636 12637 13700
rect 12571 13635 12637 13636
rect 4868 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5188 13088
rect 4868 12000 5188 13024
rect 4868 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5188 12000
rect 4868 10912 5188 11936
rect 12755 11932 12821 11933
rect 12755 11868 12756 11932
rect 12820 11868 12821 11932
rect 12755 11867 12821 11868
rect 4868 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5188 10912
rect 4868 9824 5188 10848
rect 4868 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5188 9824
rect 4868 8736 5188 9760
rect 12758 9485 12818 11867
rect 12755 9484 12821 9485
rect 12755 9420 12756 9484
rect 12820 9420 12821 9484
rect 12755 9419 12821 9420
rect 4868 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5188 8736
rect 4868 7648 5188 8672
rect 4868 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5188 7648
rect 4868 6560 5188 7584
rect 12758 6765 12818 9419
rect 19198 8125 19258 16491
rect 23979 15468 24045 15469
rect 23979 15404 23980 15468
rect 24044 15404 24045 15468
rect 23979 15403 24045 15404
rect 20483 15332 20549 15333
rect 20483 15268 20484 15332
rect 20548 15268 20549 15332
rect 20483 15267 20549 15268
rect 19195 8124 19261 8125
rect 19195 8060 19196 8124
rect 19260 8060 19261 8124
rect 19195 8059 19261 8060
rect 12755 6764 12821 6765
rect 12755 6700 12756 6764
rect 12820 6700 12821 6764
rect 12755 6699 12821 6700
rect 4868 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5188 6560
rect 4868 5472 5188 6496
rect 4868 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5188 5472
rect 4868 4384 5188 5408
rect 20486 4861 20546 15267
rect 23982 9485 24042 15403
rect 24531 13292 24597 13293
rect 24531 13228 24532 13292
rect 24596 13228 24597 13292
rect 24531 13227 24597 13228
rect 24534 9621 24594 13227
rect 24531 9620 24597 9621
rect 24531 9556 24532 9620
rect 24596 9556 24597 9620
rect 24531 9555 24597 9556
rect 23979 9484 24045 9485
rect 23979 9420 23980 9484
rect 24044 9420 24045 9484
rect 23979 9419 24045 9420
rect 20483 4860 20549 4861
rect 20483 4796 20484 4860
rect 20548 4796 20549 4860
rect 20483 4795 20549 4796
rect 4868 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5188 4384
rect 4868 3296 5188 4320
rect 4868 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5188 3296
rect 4868 2208 5188 3232
rect 4868 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5188 2208
rect 4868 2128 5188 2144
use sky130_fd_sc_hd__inv_2  _0621_
timestamp 1
transform 1 0 20884 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0622_
timestamp 1
transform -1 0 24656 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0623_
timestamp 1
transform -1 0 13432 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0624_
timestamp 1
transform 1 0 11132 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0625_
timestamp 1
transform -1 0 7176 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0626_
timestamp 1
transform 1 0 5244 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0627_
timestamp 1
transform 1 0 4416 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0628_
timestamp 1
transform 1 0 4232 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0629_
timestamp 1
transform 1 0 7636 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0630_
timestamp 1
transform 1 0 3220 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0631_
timestamp 1
transform 1 0 10120 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0632_
timestamp 1
transform 1 0 5520 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0633_
timestamp 1
transform 1 0 11592 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0634_
timestamp 1
transform 1 0 15824 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0635_
timestamp 1
transform 1 0 15180 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0636_
timestamp 1
transform 1 0 12788 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0637_
timestamp 1
transform 1 0 13340 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0638_
timestamp 1
transform -1 0 16560 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0639_
timestamp 1
transform 1 0 18584 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0640_
timestamp 1
transform -1 0 20608 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0641_
timestamp 1
transform 1 0 24104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0642_
timestamp 1
transform -1 0 20056 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0643_
timestamp 1
transform -1 0 22632 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0644_
timestamp 1
transform -1 0 23552 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0645_
timestamp 1
transform -1 0 24380 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0646_
timestamp 1
transform -1 0 21252 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0647_
timestamp 1
transform -1 0 21712 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0648_
timestamp 1
transform 1 0 22448 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0649_
timestamp 1
transform 1 0 18952 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0650_
timestamp 1
transform -1 0 18216 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0651_
timestamp 1
transform -1 0 16836 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0652_
timestamp 1
transform 1 0 15088 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0653_
timestamp 1
transform 1 0 13708 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0654_
timestamp 1
transform 1 0 13248 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0655_
timestamp 1
transform 1 0 13708 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0656_
timestamp 1
transform -1 0 13616 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0657_
timestamp 1
transform 1 0 16284 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0658_
timestamp 1
transform -1 0 25024 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0659_
timestamp 1
transform -1 0 23460 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _0660_
timestamp 1
transform -1 0 23184 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0661_
timestamp 1
transform -1 0 22724 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_2  _0662_
timestamp 1
transform -1 0 27048 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0663_
timestamp 1
transform -1 0 26588 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0664_
timestamp 1
transform -1 0 26036 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0665_
timestamp 1
transform -1 0 26128 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0666_
timestamp 1
transform 1 0 24656 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0667_
timestamp 1
transform 1 0 25024 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _0668_
timestamp 1
transform -1 0 26588 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_1  _0669_
timestamp 1
transform 1 0 25208 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0670_
timestamp 1
transform -1 0 26036 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _0671_
timestamp 1
transform 1 0 25576 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0672_
timestamp 1
transform -1 0 20516 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0673_
timestamp 1
transform -1 0 20884 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a41o_1  _0674_
timestamp 1
transform 1 0 24932 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _0675_
timestamp 1
transform -1 0 25484 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0676_
timestamp 1
transform -1 0 24288 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _0677_
timestamp 1
transform -1 0 13524 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0678_
timestamp 1
transform 1 0 4876 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _0679_
timestamp 1
transform 1 0 1656 0 1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _0680_
timestamp 1
transform 1 0 2852 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _0681_
timestamp 1
transform 1 0 1656 0 1 26112
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _0682_
timestamp 1
transform 1 0 2300 0 1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _0683_
timestamp 1
transform -1 0 3680 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0684_
timestamp 1
transform -1 0 4508 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _0685_
timestamp 1
transform 1 0 3772 0 1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__a31o_1  _0686_
timestamp 1
transform -1 0 4692 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0687_
timestamp 1
transform 1 0 5336 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0688_
timestamp 1
transform 1 0 2024 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0689_
timestamp 1
transform -1 0 3220 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0690_
timestamp 1
transform 1 0 2760 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0691_
timestamp 1
transform -1 0 4048 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0692_
timestamp 1
transform 1 0 3772 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0693_
timestamp 1
transform 1 0 4968 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0694_
timestamp 1
transform 1 0 5060 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _0695_
timestamp 1
transform 1 0 5152 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__o21bai_1  _0696_
timestamp 1
transform 1 0 3220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0697_
timestamp 1
transform 1 0 4968 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0698_
timestamp 1
transform -1 0 6348 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0699_
timestamp 1
transform -1 0 6072 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0700_
timestamp 1
transform -1 0 5612 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0701_
timestamp 1
transform 1 0 4508 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0702_
timestamp 1
transform -1 0 6256 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0703_
timestamp 1
transform -1 0 5336 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0704_
timestamp 1
transform 1 0 5612 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0705_
timestamp 1
transform -1 0 6716 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _0706_
timestamp 1
transform 1 0 6072 0 1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _0707_
timestamp 1
transform 1 0 7268 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0708_
timestamp 1
transform -1 0 5796 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0709_
timestamp 1
transform 1 0 6624 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0710_
timestamp 1
transform 1 0 5980 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0711_
timestamp 1
transform 1 0 6900 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0712_
timestamp 1
transform 1 0 6256 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0713_
timestamp 1
transform 1 0 7176 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0714_
timestamp 1
transform 1 0 7268 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0715_
timestamp 1
transform -1 0 8280 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0716_
timestamp 1
transform 1 0 9108 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0717_
timestamp 1
transform 1 0 7728 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0718_
timestamp 1
transform 1 0 8648 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0719_
timestamp 1
transform 1 0 5428 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0720_
timestamp 1
transform 1 0 1656 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0721_
timestamp 1
transform 1 0 3128 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0722_
timestamp 1
transform -1 0 9936 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0723_
timestamp 1
transform -1 0 4416 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0724_
timestamp 1
transform 1 0 1656 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0725_
timestamp 1
transform -1 0 2484 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0726_
timestamp 1
transform 1 0 2300 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0727_
timestamp 1
transform 1 0 2944 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0728_
timestamp 1
transform -1 0 4692 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0729_
timestamp 1
transform 1 0 2484 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0730_
timestamp 1
transform -1 0 4416 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0731_
timestamp 1
transform -1 0 3588 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0732_
timestamp 1
transform 1 0 4876 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0733_
timestamp 1
transform 1 0 1656 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0734_
timestamp 1
transform 1 0 2300 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0735_
timestamp 1
transform 1 0 1656 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0736_
timestamp 1
transform 1 0 3680 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0737_
timestamp 1
transform 1 0 2024 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0738_
timestamp 1
transform 1 0 2668 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0739_
timestamp 1
transform 1 0 4324 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0740_
timestamp 1
transform 1 0 3680 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o31ai_2  _0741_
timestamp 1
transform -1 0 5520 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__a31o_1  _0742_
timestamp 1
transform 1 0 2760 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0743_
timestamp 1
transform 1 0 2760 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0744_
timestamp 1
transform -1 0 4692 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _0745_
timestamp 1
transform -1 0 2852 0 -1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _0746_
timestamp 1
transform 1 0 2024 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _0747_
timestamp 1
transform 1 0 1656 0 -1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _0748_
timestamp 1
transform -1 0 3404 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _0749_
timestamp 1
transform 1 0 1932 0 -1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _0750_
timestamp 1
transform 1 0 2300 0 1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _0751_
timestamp 1
transform 1 0 3404 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _0752_
timestamp 1
transform 1 0 2484 0 1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _0753_
timestamp 1
transform 1 0 4140 0 1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _0754_
timestamp 1
transform 1 0 6348 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _0755_
timestamp 1
transform 1 0 5060 0 -1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _0756_
timestamp 1
transform 1 0 6072 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _0757_
timestamp 1
transform -1 0 4416 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0758_
timestamp 1
transform 1 0 3404 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0759_
timestamp 1
transform 1 0 4784 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _0760_
timestamp 1
transform -1 0 2852 0 -1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _0761_
timestamp 1
transform 1 0 2208 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _0762_
timestamp 1
transform 1 0 1748 0 1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _0763_
timestamp 1
transform -1 0 3128 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _0764_
timestamp 1
transform 1 0 2300 0 1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _0765_
timestamp 1
transform 1 0 3036 0 -1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__a31o_1  _0766_
timestamp 1
transform -1 0 3496 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0767_
timestamp 1
transform 1 0 3772 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _0768_
timestamp 1
transform 1 0 3772 0 1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_1  _0769_
timestamp 1
transform 1 0 4232 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0770_
timestamp 1
transform 1 0 5428 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_2  _0771_
timestamp 1
transform 1 0 4968 0 1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_1  _0772_
timestamp 1
transform 1 0 5612 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0773_
timestamp 1
transform 1 0 6900 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0774_
timestamp 1
transform -1 0 6256 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0775_
timestamp 1
transform -1 0 5520 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0776_
timestamp 1
transform -1 0 4876 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0777_
timestamp 1
transform 1 0 2576 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0778_
timestamp 1
transform 1 0 4324 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0779_
timestamp 1
transform -1 0 6624 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0780_
timestamp 1
transform 1 0 4600 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0781_
timestamp 1
transform 1 0 5244 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0782_
timestamp 1
transform 1 0 3772 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0783_
timestamp 1
transform 1 0 5152 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0784_
timestamp 1
transform 1 0 4876 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _0785_
timestamp 1
transform -1 0 6348 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0786_
timestamp 1
transform 1 0 4784 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_1  _0787_
timestamp 1
transform -1 0 6256 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0788_
timestamp 1
transform 1 0 6348 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a21boi_2  _0789_
timestamp 1
transform 1 0 6900 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_2  _0790_
timestamp 1
transform 1 0 6348 0 1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _0791_
timestamp 1
transform -1 0 7452 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _0792_
timestamp 1
transform 1 0 7452 0 -1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_1  _0793_
timestamp 1
transform 1 0 7176 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0794_
timestamp 1
transform 1 0 5520 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0795_
timestamp 1
transform 1 0 5428 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0796_
timestamp 1
transform 1 0 8556 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0797_
timestamp 1
transform 1 0 8464 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0798_
timestamp 1
transform 1 0 8280 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0799_
timestamp 1
transform -1 0 8832 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0800_
timestamp 1
transform -1 0 10396 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0801_
timestamp 1
transform 1 0 7820 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0802_
timestamp 1
transform -1 0 8740 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _0803_
timestamp 1
transform -1 0 8556 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0804_
timestamp 1
transform 1 0 7360 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0805_
timestamp 1
transform 1 0 7912 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0806_
timestamp 1
transform 1 0 6348 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0807_
timestamp 1
transform 1 0 8096 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0808_
timestamp 1
transform 1 0 7820 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0809_
timestamp 1
transform 1 0 8924 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0810_
timestamp 1
transform 1 0 8740 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0811_
timestamp 1
transform -1 0 8280 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0812_
timestamp 1
transform 1 0 7636 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0813_
timestamp 1
transform 1 0 8464 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0814_
timestamp 1
transform 1 0 9936 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0815_
timestamp 1
transform -1 0 9844 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0816_
timestamp 1
transform -1 0 9660 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0817_
timestamp 1
transform -1 0 10028 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_2  _0818_
timestamp 1
transform -1 0 9568 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0819_
timestamp 1
transform 1 0 9200 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_2  _0820_
timestamp 1
transform -1 0 7636 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _0821_
timestamp 1
transform -1 0 8832 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _0822_
timestamp 1
transform -1 0 8832 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_4  _0823_
timestamp 1
transform 1 0 6164 0 1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__o31ai_4  _0824_
timestamp 1
transform -1 0 5428 0 -1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__a31o_1  _0825_
timestamp 1
transform -1 0 3956 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0826_
timestamp 1
transform 1 0 3772 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _0827_
timestamp 1
transform 1 0 1932 0 -1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _0828_
timestamp 1
transform -1 0 3956 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _0829_
timestamp 1
transform 1 0 2484 0 -1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _0830_
timestamp 1
transform 1 0 3312 0 -1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _0831_
timestamp 1
transform 1 0 5152 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _0832_
timestamp 1
transform 1 0 3956 0 -1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _0833_
timestamp 1
transform 1 0 4692 0 -1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _0834_
timestamp 1
transform -1 0 5336 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_4  _0835_
timestamp 1
transform 1 0 5336 0 1 16320
box -38 -48 2062 592
use sky130_fd_sc_hd__xnor2_4  _0836_
timestamp 1
transform 1 0 6440 0 -1 16320
box -38 -48 2062 592
use sky130_fd_sc_hd__or2_1  _0837_
timestamp 1
transform 1 0 8372 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_4  _0838_
timestamp 1
transform 1 0 7912 0 -1 15232
box -38 -48 2062 592
use sky130_fd_sc_hd__o31ai_4  _0839_
timestamp 1
transform 1 0 4232 0 1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__a31o_1  _0840_
timestamp 1
transform -1 0 4416 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _0841_
timestamp 1
transform 1 0 3864 0 -1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _0842_
timestamp 1
transform -1 0 5060 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _0843_
timestamp 1
transform 1 0 4508 0 -1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _0844_
timestamp 1
transform 1 0 5060 0 -1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _0845_
timestamp 1
transform 1 0 6348 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_4  _0846_
timestamp 1
transform 1 0 5796 0 1 18496
box -38 -48 2062 592
use sky130_fd_sc_hd__xnor2_4  _0847_
timestamp 1
transform 1 0 6624 0 1 17408
box -38 -48 2062 592
use sky130_fd_sc_hd__a21boi_4  _0848_
timestamp 1
transform 1 0 6348 0 -1 17408
box -38 -48 1418 592
use sky130_fd_sc_hd__xnor2_4  _0849_
timestamp 1
transform 1 0 7728 0 -1 17408
box -38 -48 2062 592
use sky130_fd_sc_hd__nor2_1  _0850_
timestamp 1
transform -1 0 9384 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _0851_
timestamp 1
transform 1 0 5244 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _0852_
timestamp 1
transform 1 0 5336 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0853_
timestamp 1
transform 1 0 6900 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0854_
timestamp 1
transform 1 0 6256 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0855_
timestamp 1
transform 1 0 7360 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a21boi_2  _0856_
timestamp 1
transform 1 0 6808 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0857_
timestamp 1
transform -1 0 9200 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0858_
timestamp 1
transform 1 0 8464 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0859_
timestamp 1
transform 1 0 9660 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_2  _0860_
timestamp 1
transform 1 0 7084 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_2  _0861_
timestamp 1
transform 1 0 7084 0 -1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _0862_
timestamp 1
transform 1 0 8924 0 1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _0863_
timestamp 1
transform -1 0 10212 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0864_
timestamp 1
transform 1 0 7544 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0865_
timestamp 1
transform 1 0 7728 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0866_
timestamp 1
transform 1 0 9384 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0867_
timestamp 1
transform -1 0 8464 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0868_
timestamp 1
transform 1 0 8188 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__a41oi_4  _0869_
timestamp 1
transform 1 0 8924 0 1 17408
box -38 -48 2062 592
use sky130_fd_sc_hd__nand2_1  _0870_
timestamp 1
transform 1 0 9200 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0871_
timestamp 1
transform -1 0 10028 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _0872_
timestamp 1
transform 1 0 6992 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _0873_
timestamp 1
transform 1 0 6348 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0874_
timestamp 1
transform 1 0 7084 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__o31ai_1  _0875_
timestamp 1
transform 1 0 6532 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0876_
timestamp 1
transform 1 0 7452 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0877_
timestamp 1
transform 1 0 7728 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0878_
timestamp 1
transform 1 0 7544 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0879_
timestamp 1
transform 1 0 8004 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _0880_
timestamp 1
transform -1 0 8648 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__nor3b_1  _0881_
timestamp 1
transform -1 0 9200 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0882_
timestamp 1
transform 1 0 8924 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _0883_
timestamp 1
transform -1 0 11316 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0884_
timestamp 1
transform 1 0 9476 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _0885_
timestamp 1
transform -1 0 11960 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nand4_2  _0886_
timestamp 1
transform 1 0 10580 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__a31o_1  _0887_
timestamp 1
transform 1 0 10488 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _0888_
timestamp 1
transform 1 0 9936 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0889_
timestamp 1
transform -1 0 11960 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _0890_
timestamp 1
transform 1 0 10304 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _0891_
timestamp 1
transform 1 0 10672 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _0892_
timestamp 1
transform -1 0 10304 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__nand3_1  _0893_
timestamp 1
transform 1 0 9752 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0894_
timestamp 1
transform 1 0 10120 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0895_
timestamp 1
transform 1 0 10396 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0896_
timestamp 1
transform -1 0 9384 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0897_
timestamp 1
transform -1 0 9476 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _0898_
timestamp 1
transform -1 0 8832 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0899_
timestamp 1
transform 1 0 9292 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0900_
timestamp 1
transform 1 0 9844 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0901_
timestamp 1
transform 1 0 9384 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _0902_
timestamp 1
transform -1 0 10488 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0903_
timestamp 1
transform -1 0 9108 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0904_
timestamp 1
transform 1 0 9476 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _0905_
timestamp 1
transform 1 0 10028 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0906_
timestamp 1
transform -1 0 11040 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0907_
timestamp 1
transform 1 0 12604 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0908_
timestamp 1
transform 1 0 12512 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0909_
timestamp 1
transform 1 0 11960 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0910_
timestamp 1
transform -1 0 12788 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0911_
timestamp 1
transform 1 0 12052 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_2  _0912_
timestamp 1
transform 1 0 11592 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0913_
timestamp 1
transform -1 0 12880 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0914_
timestamp 1
transform 1 0 12236 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__o211ai_4  _0915_
timestamp 1
transform 1 0 12236 0 1 23936
box -38 -48 1602 592
use sky130_fd_sc_hd__o21a_1  _0916_
timestamp 1
transform -1 0 13432 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0917_
timestamp 1
transform 1 0 14812 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0918_
timestamp 1
transform 1 0 14352 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0919_
timestamp 1
transform -1 0 14628 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0920_
timestamp 1
transform 1 0 14904 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_2  _0921_
timestamp 1
transform 1 0 14812 0 -1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__a211o_1  _0922_
timestamp 1
transform -1 0 12972 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0923_
timestamp 1
transform -1 0 12328 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0924_
timestamp 1
transform 1 0 12880 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0925_
timestamp 1
transform -1 0 12880 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0926_
timestamp 1
transform 1 0 11776 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0927_
timestamp 1
transform -1 0 13248 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0928_
timestamp 1
transform 1 0 13064 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0929_
timestamp 1
transform 1 0 14076 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nor3b_1  _0930_
timestamp 1
transform -1 0 16560 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _0931_
timestamp 1
transform 1 0 16376 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0932_
timestamp 1
transform -1 0 10028 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _0933_
timestamp 1
transform 1 0 15548 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0934_
timestamp 1
transform -1 0 15548 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__nand3b_1  _0935_
timestamp 1
transform 1 0 15824 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _0936_
timestamp 1
transform 1 0 15088 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0937_
timestamp 1
transform 1 0 15732 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0938_
timestamp 1
transform -1 0 17204 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0939_
timestamp 1
transform 1 0 17204 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0940_
timestamp 1
transform 1 0 16284 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o211ai_1  _0941_
timestamp 1
transform 1 0 10028 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0942_
timestamp 1
transform 1 0 14076 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0943_
timestamp 1
transform -1 0 18492 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0944_
timestamp 1
transform 1 0 17756 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0945_
timestamp 1
transform -1 0 11040 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _0946_
timestamp 1
transform 1 0 10028 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0947_
timestamp 1
transform 1 0 18492 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0948_
timestamp 1
transform -1 0 20424 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _0949_
timestamp 1
transform 1 0 18768 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_2  _0950_
timestamp 1
transform 1 0 9476 0 1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _0951_
timestamp 1
transform 1 0 21252 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0952_
timestamp 1
transform 1 0 19228 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a311oi_1  _0953_
timestamp 1
transform 1 0 16652 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a311o_1  _0954_
timestamp 1
transform 1 0 17112 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__and4bb_1  _0955_
timestamp 1
transform 1 0 16192 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__or3b_1  _0956_
timestamp 1
transform 1 0 13892 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a211oi_2  _0957_
timestamp 1
transform -1 0 15548 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _0958_
timestamp 1
transform -1 0 15180 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_4  _0959_
timestamp 1
transform -1 0 16008 0 1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__or3_1  _0960_
timestamp 1
transform 1 0 15088 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0961_
timestamp 1
transform -1 0 21252 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0962_
timestamp 1
transform -1 0 20700 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _0963_
timestamp 1
transform -1 0 20056 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nand4_1  _0964_
timestamp 1
transform -1 0 17756 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0965_
timestamp 1
transform -1 0 9660 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0966_
timestamp 1
transform 1 0 10948 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_2  _0967_
timestamp 1
transform 1 0 9844 0 -1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _0968_
timestamp 1
transform -1 0 18952 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _0969_
timestamp 1
transform 1 0 9752 0 -1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_1  _0970_
timestamp 1
transform -1 0 21528 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0971_
timestamp 1
transform 1 0 20424 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0972_
timestamp 1
transform 1 0 20792 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_2  _0973_
timestamp 1
transform -1 0 9292 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_4  _0974_
timestamp 1
transform 1 0 9292 0 -1 16320
box -38 -48 2062 592
use sky130_fd_sc_hd__inv_2  _0975_
timestamp 1
transform 1 0 16652 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0976_
timestamp 1
transform 1 0 21252 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0977_
timestamp 1
transform -1 0 21988 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_4  _0978_
timestamp 1
transform 1 0 9200 0 1 15232
box -38 -48 2062 592
use sky130_fd_sc_hd__xnor2_1  _0979_
timestamp 1
transform -1 0 21436 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _0980_
timestamp 1
transform -1 0 21068 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _0981_
timestamp 1
transform 1 0 8648 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_2  _0982_
timestamp 1
transform 1 0 8924 0 1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _0983_
timestamp 1
transform -1 0 19596 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0984_
timestamp 1
transform 1 0 20700 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0985_
timestamp 1
transform 1 0 20976 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _0986_
timestamp 1
transform 1 0 8924 0 -1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _0987_
timestamp 1
transform -1 0 18860 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0988_
timestamp 1
transform 1 0 19320 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _0989_
timestamp 1
transform -1 0 20608 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0990_
timestamp 1
transform 1 0 9016 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _0991_
timestamp 1
transform 1 0 10396 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0992_
timestamp 1
transform -1 0 17112 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0993_
timestamp 1
transform 1 0 9476 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0994_
timestamp 1
transform 1 0 9936 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0995_
timestamp 1
transform -1 0 16560 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0996_
timestamp 1
transform 1 0 9016 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0997_
timestamp 1
transform 1 0 9476 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0998_
timestamp 1
transform 1 0 14628 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0999_
timestamp 1
transform 1 0 15640 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1000_
timestamp 1
transform 1 0 8740 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1001_
timestamp 1
transform 1 0 9384 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1002_
timestamp 1
transform 1 0 13800 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1003_
timestamp 1
transform -1 0 14168 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1004_
timestamp 1
transform -1 0 12880 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1005_
timestamp 1
transform 1 0 13064 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1006_
timestamp 1
transform -1 0 13800 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1007_
timestamp 1
transform 1 0 11592 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1008_
timestamp 1
transform -1 0 11776 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1009_
timestamp 1
transform -1 0 12420 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1010_
timestamp 1
transform 1 0 12052 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1011_
timestamp 1
transform 1 0 12604 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__o21ba_1  _1012_
timestamp 1
transform -1 0 14720 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1013_
timestamp 1
transform 1 0 16652 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1014_
timestamp 1
transform 1 0 8740 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _1015_
timestamp 1
transform 1 0 9568 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1016_
timestamp 1
transform 1 0 20148 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1017_
timestamp 1
transform -1 0 19964 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1018_
timestamp 1
transform -1 0 19688 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1019_
timestamp 1
transform 1 0 9292 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _1020_
timestamp 1
transform 1 0 9568 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1021_
timestamp 1
transform 1 0 17940 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o2111ai_1  _1022_
timestamp 1
transform -1 0 18952 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1023_
timestamp 1
transform 1 0 18308 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_1  _1024_
timestamp 1
transform 1 0 18676 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1025_
timestamp 1
transform -1 0 19872 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o311a_1  _1026_
timestamp 1
transform 1 0 19228 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1027_
timestamp 1
transform 1 0 20608 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1028_
timestamp 1
transform -1 0 21620 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _1029_
timestamp 1
transform 1 0 21068 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1030_
timestamp 1
transform 1 0 20608 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_2  _1031_
timestamp 1
transform 1 0 19228 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a41oi_4  _1032_
timestamp 1
transform 1 0 17112 0 -1 21760
box -38 -48 2062 592
use sky130_fd_sc_hd__a41o_1  _1033_
timestamp 1
transform 1 0 17112 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  _1034_
timestamp 1
transform -1 0 23276 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _1035_
timestamp 1
transform 1 0 23736 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1036_
timestamp 1
transform -1 0 24932 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _1037_
timestamp 1
transform 1 0 14168 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _1038_
timestamp 1
transform 1 0 14076 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1039_
timestamp 1
transform 1 0 15088 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1040_
timestamp 1
transform 1 0 17480 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1041_
timestamp 1
transform 1 0 18400 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_1  _1042_
timestamp 1
transform -1 0 18584 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_4  _1043_
timestamp 1
transform -1 0 23644 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__and4_1  _1044_
timestamp 1
transform 1 0 9292 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1045_
timestamp 1
transform -1 0 10948 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1046_
timestamp 1
transform 1 0 10948 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1047_
timestamp 1
transform 1 0 19688 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1048_
timestamp 1
transform 1 0 22264 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_2  _1049_
timestamp 1
transform 1 0 23644 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1050_
timestamp 1
transform -1 0 22448 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1051_
timestamp 1
transform -1 0 23552 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__o311a_1  _1052_
timestamp 1
transform -1 0 24288 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1053_
timestamp 1
transform 1 0 24748 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1054_
timestamp 1
transform -1 0 24656 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1055_
timestamp 1
transform 1 0 24288 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o21bai_1  _1056_
timestamp 1
transform -1 0 24564 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1057_
timestamp 1
transform -1 0 25392 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _1058_
timestamp 1
transform 1 0 23000 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1059_
timestamp 1
transform 1 0 24012 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1060_
timestamp 1
transform 1 0 22908 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1061_
timestamp 1
transform 1 0 23184 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1062_
timestamp 1
transform -1 0 23184 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1063_
timestamp 1
transform -1 0 24288 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1064_
timestamp 1
transform 1 0 24380 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1065_
timestamp 1
transform -1 0 24288 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _1066_
timestamp 1
transform 1 0 21896 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1067_
timestamp 1
transform 1 0 22448 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1068_
timestamp 1
transform 1 0 23644 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1069_
timestamp 1
transform 1 0 21344 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1070_
timestamp 1
transform 1 0 22908 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1071_
timestamp 1
transform 1 0 22448 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1072_
timestamp 1
transform 1 0 24840 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1073_
timestamp 1
transform 1 0 15640 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1074_
timestamp 1
transform 1 0 14076 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1075_
timestamp 1
transform 1 0 14812 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1076_
timestamp 1
transform 1 0 15272 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a31oi_1  _1077_
timestamp 1
transform 1 0 14444 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1078_
timestamp 1
transform 1 0 12420 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1079_
timestamp 1
transform -1 0 13800 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1080_
timestamp 1
transform 1 0 13616 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__o41a_1  _1081_
timestamp 1
transform 1 0 12696 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _1082_
timestamp 1
transform 1 0 13064 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1083_
timestamp 1
transform 1 0 11868 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _1084_
timestamp 1
transform 1 0 11960 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1085_
timestamp 1
transform -1 0 13708 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1086_
timestamp 1
transform 1 0 13432 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o41a_1  _1087_
timestamp 1
transform 1 0 12604 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _1088_
timestamp 1
transform 1 0 12236 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1089_
timestamp 1
transform 1 0 11868 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1090_
timestamp 1
transform 1 0 12420 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1091_
timestamp 1
transform 1 0 12512 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1092_
timestamp 1
transform 1 0 12788 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1093_
timestamp 1
transform -1 0 12052 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1094_
timestamp 1
transform -1 0 13248 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1095_
timestamp 1
transform 1 0 13156 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1096_
timestamp 1
transform 1 0 12328 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1097_
timestamp 1
transform -1 0 11224 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1098_
timestamp 1
transform 1 0 13064 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1099_
timestamp 1
transform 1 0 12972 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1100_
timestamp 1
transform -1 0 13064 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__o41a_1  _1101_
timestamp 1
transform 1 0 13432 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__a221oi_2  _1102_
timestamp 1
transform 1 0 12144 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_1  _1103_
timestamp 1
transform 1 0 15364 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1104_
timestamp 1
transform -1 0 14904 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1105_
timestamp 1
transform 1 0 16284 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1106_
timestamp 1
transform -1 0 16284 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _1107_
timestamp 1
transform 1 0 14904 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1108_
timestamp 1
transform -1 0 14536 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1109_
timestamp 1
transform -1 0 18676 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1110_
timestamp 1
transform 1 0 15364 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1111_
timestamp 1
transform -1 0 15640 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1112_
timestamp 1
transform 1 0 15824 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1113_
timestamp 1
transform 1 0 16008 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a31oi_1  _1114_
timestamp 1
transform 1 0 15272 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1115_
timestamp 1
transform 1 0 17296 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1116_
timestamp 1
transform 1 0 16652 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1117_
timestamp 1
transform -1 0 17480 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _1118_
timestamp 1
transform -1 0 17388 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1119_
timestamp 1
transform 1 0 17940 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a31oi_1  _1120_
timestamp 1
transform 1 0 16744 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1121_
timestamp 1
transform -1 0 19136 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1122_
timestamp 1
transform 1 0 19412 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1123_
timestamp 1
transform 1 0 19872 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o41a_1  _1124_
timestamp 1
transform 1 0 19228 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__a221oi_4  _1125_
timestamp 1
transform 1 0 18216 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__a211o_1  _1126_
timestamp 1
transform -1 0 21344 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1127_
timestamp 1
transform 1 0 20700 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _1128_
timestamp 1
transform 1 0 21804 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1129_
timestamp 1
transform -1 0 20700 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1130_
timestamp 1
transform 1 0 21344 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _1131_
timestamp 1
transform 1 0 20976 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1132_
timestamp 1
transform 1 0 20884 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1133_
timestamp 1
transform -1 0 20516 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o41a_1  _1134_
timestamp 1
transform 1 0 21804 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _1135_
timestamp 1
transform 1 0 20884 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1136_
timestamp 1
transform 1 0 20424 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1137_
timestamp 1
transform 1 0 20148 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1138_
timestamp 1
transform 1 0 21804 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1139_
timestamp 1
transform 1 0 21528 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1140_
timestamp 1
transform -1 0 21712 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1141_
timestamp 1
transform -1 0 20976 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _1142_
timestamp 1
transform 1 0 19596 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1143_
timestamp 1
transform -1 0 19688 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1144_
timestamp 1
transform -1 0 22816 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1145_
timestamp 1
transform 1 0 24380 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _1146_
timestamp 1
transform 1 0 24380 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a221oi_2  _1147_
timestamp 1
transform -1 0 23920 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__a211o_1  _1148_
timestamp 1
transform 1 0 22448 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1149_
timestamp 1
transform -1 0 24840 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1150_
timestamp 1
transform 1 0 24840 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__o41a_1  _1151_
timestamp 1
transform 1 0 23460 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _1152_
timestamp 1
transform -1 0 24196 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1153_
timestamp 1
transform 1 0 23092 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1154_
timestamp 1
transform 1 0 22080 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1155_
timestamp 1
transform -1 0 24932 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1156_
timestamp 1
transform 1 0 24380 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1157_
timestamp 1
transform -1 0 24472 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1158_
timestamp 1
transform 1 0 23184 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__a211oi_2  _1159_
timestamp 1
transform -1 0 24288 0 1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__xnor2_1  _1160_
timestamp 1
transform -1 0 23276 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _1161_
timestamp 1
transform -1 0 18952 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _1162_
timestamp 1
transform 1 0 18124 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1163_
timestamp 1
transform 1 0 17848 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1164_
timestamp 1
transform 1 0 21896 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1165_
timestamp 1
transform -1 0 24104 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1166_
timestamp 1
transform -1 0 23644 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _1167_
timestamp 1
transform -1 0 23644 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1168_
timestamp 1
transform 1 0 21804 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1169_
timestamp 1
transform 1 0 22540 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1170_
timestamp 1
transform -1 0 22540 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1171_
timestamp 1
transform -1 0 21252 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1172_
timestamp 1
transform -1 0 21528 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1173_
timestamp 1
transform -1 0 20792 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o221ai_2  _1174_
timestamp 1
transform -1 0 20608 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__a21oi_1  _1175_
timestamp 1
transform 1 0 21068 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1176_
timestamp 1
transform -1 0 20332 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1177_
timestamp 1
transform 1 0 18584 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1178_
timestamp 1
transform 1 0 19136 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _1179_
timestamp 1
transform 1 0 19228 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1180_
timestamp 1
transform 1 0 18400 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1181_
timestamp 1
transform -1 0 18952 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1182_
timestamp 1
transform 1 0 18860 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1183_
timestamp 1
transform 1 0 16744 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1184_
timestamp 1
transform 1 0 17204 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1185_
timestamp 1
transform 1 0 17112 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o221ai_4  _1186_
timestamp 1
transform -1 0 18584 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__a21oi_1  _1187_
timestamp 1
transform -1 0 16652 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1188_
timestamp 1
transform -1 0 16468 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1189_
timestamp 1
transform 1 0 12972 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1190_
timestamp 1
transform 1 0 13432 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1191_
timestamp 1
transform -1 0 12880 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1192_
timestamp 1
transform -1 0 13432 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1193_
timestamp 1
transform 1 0 14076 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1194_
timestamp 1
transform 1 0 12788 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1195_
timestamp 1
transform -1 0 11776 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1196_
timestamp 1
transform -1 0 14260 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1197_
timestamp 1
transform -1 0 13892 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1198_
timestamp 1
transform -1 0 13616 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a41oi_1  _1199_
timestamp 1
transform -1 0 13156 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a221oi_2  _1200_
timestamp 1
transform 1 0 11776 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__xnor2_1  _1201_
timestamp 1
transform 1 0 13340 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _1202_
timestamp 1
transform -1 0 15916 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1203_
timestamp 1
transform -1 0 16008 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  _1204_
timestamp 1
transform -1 0 14996 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a211oi_1  _1205_
timestamp 1
transform -1 0 12236 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1206_
timestamp 1
transform 1 0 13156 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1207_
timestamp 1
transform 1 0 12880 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a41o_1  _1208_
timestamp 1
transform 1 0 12604 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1209_
timestamp 1
transform 1 0 12696 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1210_
timestamp 1
transform -1 0 24012 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1211_
timestamp 1
transform -1 0 19320 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1212_
timestamp 1
transform 1 0 22632 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a311o_1  _1213_
timestamp 1
transform 1 0 23644 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_1  _1214_
timestamp 1
transform 1 0 22908 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1215_
timestamp 1
transform 1 0 16836 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o22ai_1  _1216_
timestamp 1
transform -1 0 16192 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_1  _1217_
timestamp 1
transform -1 0 17940 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _1218_
timestamp 1
transform -1 0 12236 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1219_
timestamp 1
transform 1 0 16744 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1220_
timestamp 1
transform -1 0 21896 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1221_
timestamp 1
transform -1 0 21620 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1222_
timestamp 1
transform -1 0 19780 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__o2111ai_1  _1223_
timestamp 1
transform 1 0 20240 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _1224_
timestamp 1
transform -1 0 16560 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1225_
timestamp 1
transform 1 0 13432 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1226_
timestamp 1
transform -1 0 15640 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a2111o_1  _1227_
timestamp 1
transform 1 0 15364 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _1228_
timestamp 1
transform 1 0 20056 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1229_
timestamp 1
transform 1 0 18400 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1230_
timestamp 1
transform 1 0 13064 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1231_
timestamp 1
transform -1 0 17572 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__o2111ai_1  _1232_
timestamp 1
transform -1 0 17296 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a311o_1  _1233_
timestamp 1
transform 1 0 15732 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a311o_1  _1234_
timestamp 1
transform -1 0 22264 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1235_
timestamp 1
transform -1 0 13248 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o2111ai_1  _1236_
timestamp 1
transform 1 0 15088 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1237_
timestamp 1
transform 1 0 16192 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _1238_
timestamp 1
transform -1 0 12328 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a2111o_1  _1239_
timestamp 1
transform -1 0 15364 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__a2bb2o_1  _1240_
timestamp 1
transform 1 0 12420 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1241_
timestamp 1
transform 1 0 11500 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _1242_
timestamp 1
transform 1 0 16836 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1243_
timestamp 1
transform 1 0 12052 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1244_
timestamp 1
transform 1 0 12788 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _1245_
timestamp 1
transform 1 0 20056 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o31ai_1  _1246_
timestamp 1
transform 1 0 17572 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _1247_
timestamp 1
transform 1 0 18400 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__o32ai_1  _1248_
timestamp 1
transform 1 0 18032 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a311o_1  _1249_
timestamp 1
transform 1 0 14904 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__o31ai_1  _1250_
timestamp 1
transform 1 0 14536 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1251_
timestamp 1
transform -1 0 18216 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1252_
timestamp 1
transform 1 0 16928 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1253_
timestamp 1
transform -1 0 22080 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  _1254_
timestamp 1
transform -1 0 25576 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _1255_
timestamp 1
transform -1 0 26128 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1256_
timestamp 1
transform 1 0 22816 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1257_
timestamp 1
transform -1 0 26772 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1258_
timestamp 1
transform 1 0 26772 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_1  _1259_
timestamp 1
transform 1 0 26128 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1260_
timestamp 1
transform -1 0 27232 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_1  _1261_
timestamp 1
transform -1 0 19596 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1262_
timestamp 1
transform 1 0 25668 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1263_
timestamp 1
transform 1 0 26956 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _1264_
timestamp 1
transform -1 0 26404 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1265_
timestamp 1
transform -1 0 18768 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1266_
timestamp 1
transform -1 0 18860 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_1  _1267_
timestamp 1
transform 1 0 26036 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1268_
timestamp 1
transform -1 0 27324 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1269_
timestamp 1
transform -1 0 20056 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_1  _1270_
timestamp 1
transform -1 0 17940 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1271_
timestamp 1
transform 1 0 17204 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _1272_
timestamp 1
transform -1 0 21528 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _1273_
timestamp 1
transform 1 0 20516 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1274_
timestamp 1
transform -1 0 20332 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1275_
timestamp 1
transform -1 0 18584 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1276_
timestamp 1
transform -1 0 22264 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_1  _1277_
timestamp 1
transform 1 0 24104 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1278_
timestamp 1
transform -1 0 24288 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_1  _1279_
timestamp 1
transform -1 0 20332 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1280_
timestamp 1
transform 1 0 20332 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__or4bb_1  _1281_
timestamp 1
transform 1 0 25208 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1282_
timestamp 1
transform 1 0 26128 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__o311a_1  _1283_
timestamp 1
transform -1 0 21068 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__and4b_1  _1284_
timestamp 1
transform 1 0 23092 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__or4bb_1  _1285_
timestamp 1
transform 1 0 24380 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1286_
timestamp 1
transform 1 0 25300 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1287_
timestamp 1
transform -1 0 19044 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _1288_
timestamp 1
transform -1 0 19872 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1289_
timestamp 1
transform -1 0 20056 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__and4bb_1  _1290_
timestamp 1
transform -1 0 22356 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__and4b_1  _1291_
timestamp 1
transform -1 0 23092 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_2  _1292_
timestamp 1
transform -1 0 26864 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1293_
timestamp 1
transform -1 0 21712 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1294_
timestamp 1
transform 1 0 21804 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1295_
timestamp 1
transform 1 0 17296 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1296_
timestamp 1
transform 1 0 26772 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1297_
timestamp 1
transform 1 0 16928 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1298_
timestamp 1
transform -1 0 21436 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1299_
timestamp 1
transform -1 0 20516 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1300_
timestamp 1
transform -1 0 25116 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1301_
timestamp 1
transform 1 0 17848 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1302_
timestamp 1
transform 1 0 25852 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_1  _1303_
timestamp 1
transform 1 0 25116 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1304_
timestamp 1
transform 1 0 26220 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1305_
timestamp 1
transform 1 0 24840 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1306_
timestamp 1
transform -1 0 18584 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _1307_
timestamp 1
transform -1 0 19596 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1308_
timestamp 1
transform 1 0 25576 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1309_
timestamp 1
transform 1 0 27048 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _1310_
timestamp 1
transform 1 0 26588 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1311_
timestamp 1
transform 1 0 26956 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__dfrtp_1  _1312_
timestamp 1
transform 1 0 22816 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1313_
timestamp 1
transform 1 0 24380 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1314_
timestamp 1
transform 1 0 25024 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1315_
timestamp 1
transform 1 0 23644 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1316_
timestamp 1
transform 1 0 23460 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1317_
timestamp 1
transform -1 0 16376 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1318_
timestamp 1
transform 1 0 11500 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1319_
timestamp 1
transform -1 0 12604 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1320_
timestamp 1
transform 1 0 11500 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1321_
timestamp 1
transform 1 0 11224 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1322_
timestamp 1
transform 1 0 14352 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1323_
timestamp 1
transform 1 0 16284 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1324_
timestamp 1
transform 1 0 16836 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1325_
timestamp 1
transform 1 0 17296 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1326_
timestamp 1
transform 1 0 20056 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1327_
timestamp 1
transform 1 0 20516 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1328_
timestamp 1
transform 1 0 19688 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1329_
timestamp 1
transform 1 0 23920 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1330_
timestamp 1
transform -1 0 26220 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1331_
timestamp 1
transform -1 0 26496 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1332_
timestamp 1
transform 1 0 17664 0 -1 17408
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1333_
timestamp 1
transform 1 0 22264 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1334_
timestamp 1
transform 1 0 19228 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1335_
timestamp 1
transform 1 0 19228 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1336_
timestamp 1
transform 1 0 15272 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1337_
timestamp 1
transform 1 0 10580 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1338_
timestamp 1
transform 1 0 10672 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1339_
timestamp 1
transform 1 0 14996 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1340_
timestamp 1
transform 1 0 12236 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1341_
timestamp 1
transform 1 0 26036 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1342_
timestamp 1
transform 1 0 25300 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1343_
timestamp 1
transform 1 0 25576 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1344_
timestamp 1
transform 1 0 22264 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1345_
timestamp 1
transform 1 0 21804 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1346_
timestamp 1
transform 1 0 21896 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1347_
timestamp 1
transform 1 0 24380 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp 1
transform -1 0 20608 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_clk
timestamp 1
transform -1 0 18860 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_clk
timestamp 1
transform 1 0 20240 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_clk
timestamp 1
transform -1 0 19136 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_clk
timestamp 1
transform 1 0 20976 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkload0
timestamp 1
transform 1 0 17020 0 -1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_2  clkload1
timestamp 1
transform 1 0 20332 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  clkload2
timestamp 1
transform 1 0 17664 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout53
timestamp 1
transform -1 0 17480 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout54
timestamp 1
transform 1 0 22908 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout55
timestamp 1
transform 1 0 16008 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout56
timestamp 1
transform 1 0 19596 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout57
timestamp 1
transform 1 0 17848 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout58
timestamp 1
transform -1 0 16928 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout59
timestamp 1
transform 1 0 13524 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout60
timestamp 1
transform -1 0 12788 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout61
timestamp 1
transform -1 0 13984 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout62
timestamp 1
transform -1 0 19228 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout63
timestamp 1
transform -1 0 20516 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout64
timestamp 1
transform -1 0 16192 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout65
timestamp 1
transform 1 0 23184 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout66
timestamp 1
transform -1 0 25852 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout67
timestamp 1
transform -1 0 23644 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout68
timestamp 1
transform -1 0 23368 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout69
timestamp 1
transform 1 0 24840 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout70
timestamp 1
transform -1 0 21252 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout71
timestamp 1
transform -1 0 26680 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout72
timestamp 1
transform -1 0 27324 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout73
timestamp 1
transform 1 0 26036 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout74
timestamp 1
transform -1 0 25760 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  fanout75
timestamp 1
transform 1 0 21988 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout76
timestamp 1
transform -1 0 23276 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout77
timestamp 1
transform -1 0 21988 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout78
timestamp 1
transform -1 0 6440 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout79
timestamp 1
transform -1 0 3220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout80
timestamp 1
transform -1 0 3680 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout81
timestamp 1
transform 1 0 12604 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout82
timestamp 1
transform -1 0 3312 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout83
timestamp 1
transform -1 0 25852 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout84
timestamp 1
transform -1 0 25116 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout85
timestamp 1
transform -1 0 25760 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout86
timestamp 1
transform -1 0 26772 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout87
timestamp 1
transform -1 0 2484 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout88
timestamp 1
transform -1 0 24196 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout89
timestamp 1
transform 1 0 22632 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout90
timestamp 1
transform 1 0 25024 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout91
timestamp 1
transform -1 0 24748 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3
timestamp 1636968456
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 1636968456
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27
timestamp 1
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1636968456
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41
timestamp 1
transform 1 0 4876 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49
timestamp 1
transform 1 0 5612 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55
timestamp 1
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1636968456
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1636968456
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91
timestamp 1636968456
transform 1 0 9476 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_103
timestamp 1
transform 1 0 10580 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111
timestamp 1
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1636968456
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 1636968456
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1636968456
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1636968456
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1636968456
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_181
timestamp 1636968456
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 1
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_197
timestamp 1636968456
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_209
timestamp 1636968456
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_221
timestamp 1
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_225
timestamp 1636968456
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_237
timestamp 1636968456
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp 1
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_253
timestamp 1636968456
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_265
timestamp 1636968456
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_277
timestamp 1
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_281
timestamp 1
transform 1 0 26956 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_289
timestamp 1
transform 1 0 27692 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1636968456
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1636968456
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1636968456
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1636968456
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 1
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1636968456
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1636968456
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1636968456
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1636968456
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1636968456
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1636968456
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1636968456
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1636968456
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1636968456
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_181
timestamp 1636968456
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_193
timestamp 1636968456
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_205
timestamp 1636968456
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp 1
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1636968456
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_237
timestamp 1636968456
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_249
timestamp 1636968456
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_261
timestamp 1636968456
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp 1
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_281
timestamp 1
transform 1 0 26956 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_289
timestamp 1
transform 1 0 27692 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1636968456
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1636968456
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1636968456
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1636968456
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1636968456
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1636968456
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1636968456
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1636968456
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1636968456
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1636968456
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1636968456
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1636968456
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1636968456
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1636968456
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1636968456
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1636968456
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_221
timestamp 1636968456
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_233
timestamp 1636968456
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 1
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1636968456
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_265
timestamp 1636968456
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_277
timestamp 1636968456
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_289
timestamp 1
transform 1 0 27692 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1636968456
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1636968456
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1636968456
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1636968456
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1636968456
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1636968456
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1636968456
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1636968456
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1636968456
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1636968456
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1636968456
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1636968456
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1636968456
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1636968456
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1636968456
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1636968456
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1636968456
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1636968456
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_249
timestamp 1636968456
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_261
timestamp 1636968456
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_281
timestamp 1
transform 1 0 26956 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_289
timestamp 1
transform 1 0 27692 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1636968456
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1636968456
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1636968456
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1636968456
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1636968456
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1636968456
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1636968456
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1636968456
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1636968456
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1636968456
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1636968456
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1636968456
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1636968456
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1636968456
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1636968456
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1636968456
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_221
timestamp 1636968456
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_233
timestamp 1636968456
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1636968456
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1636968456
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_277
timestamp 1636968456
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_289
timestamp 1
transform 1 0 27692 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1636968456
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1636968456
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1636968456
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1636968456
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1636968456
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1636968456
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1636968456
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1636968456
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1636968456
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1636968456
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1636968456
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1636968456
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1636968456
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1636968456
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1636968456
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1636968456
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1636968456
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1636968456
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_249
timestamp 1636968456
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_261
timestamp 1636968456
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_281
timestamp 1
transform 1 0 26956 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_289
timestamp 1
transform 1 0 27692 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1636968456
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1636968456
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1636968456
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1636968456
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1636968456
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1636968456
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_77
timestamp 1
transform 1 0 8188 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1636968456
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1636968456
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1636968456
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1636968456
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1636968456
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1636968456
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1636968456
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1636968456
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1636968456
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1636968456
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_221
timestamp 1636968456
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_233
timestamp 1636968456
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1636968456
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1636968456
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_277
timestamp 1
transform 1 0 26588 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_285
timestamp 1
transform 1 0 27324 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1636968456
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1636968456
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1636968456
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1636968456
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1636968456
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_69
timestamp 1
transform 1 0 7452 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_7_80
timestamp 1
transform 1 0 8464 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_90
timestamp 1636968456
transform 1 0 9384 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_102
timestamp 1
transform 1 0 10488 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_110
timestamp 1
transform 1 0 11224 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_136
timestamp 1
transform 1 0 13616 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_144
timestamp 1
transform 1 0 14352 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_166
timestamp 1
transform 1 0 16376 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_169
timestamp 1
transform 1 0 16652 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_192
timestamp 1636968456
transform 1 0 18768 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_204
timestamp 1636968456
transform 1 0 19872 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_216
timestamp 1
transform 1 0 20976 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1636968456
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1636968456
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_249
timestamp 1636968456
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_261
timestamp 1636968456
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_281
timestamp 1
transform 1 0 26956 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_287
timestamp 1
transform 1 0 27508 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1636968456
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1636968456
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1636968456
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_41
timestamp 1
transform 1 0 4876 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_8_54
timestamp 1636968456
transform 1 0 6072 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_66
timestamp 1
transform 1 0 7176 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_95
timestamp 1
transform 1 0 9844 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_101
timestamp 1636968456
transform 1 0 10396 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_113
timestamp 1
transform 1 0 11500 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_121
timestamp 1
transform 1 0 12236 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_148
timestamp 1
transform 1 0 14720 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_163
timestamp 1636968456
transform 1 0 16100 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_175
timestamp 1
transform 1 0 17204 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_197
timestamp 1
transform 1 0 19228 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_205
timestamp 1
transform 1 0 19964 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_227
timestamp 1636968456
transform 1 0 21988 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_239
timestamp 1
transform 1 0 23092 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1636968456
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1636968456
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_277
timestamp 1636968456
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_289
timestamp 1
transform 1 0 27692 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1636968456
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1636968456
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_27
timestamp 1
transform 1 0 3588 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_35
timestamp 1
transform 1 0 4324 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_60
timestamp 1636968456
transform 1 0 6624 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_72
timestamp 1
transform 1 0 7728 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_85
timestamp 1
transform 1 0 8924 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_106
timestamp 1
transform 1 0 10856 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_121
timestamp 1
transform 1 0 12236 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_125
timestamp 1
transform 1 0 12604 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_142
timestamp 1
transform 1 0 14168 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_169
timestamp 1
transform 1 0 16652 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_235
timestamp 1
transform 1 0 22724 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_239
timestamp 1
transform 1 0 23092 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_263
timestamp 1636968456
transform 1 0 25300 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_275
timestamp 1
transform 1 0 26404 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_281
timestamp 1
transform 1 0 26956 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_289
timestamp 1
transform 1 0 27692 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1636968456
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1636968456
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_29
timestamp 1
transform 1 0 3772 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_10_58
timestamp 1636968456
transform 1 0 6440 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_70
timestamp 1636968456
transform 1 0 7544 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_82
timestamp 1
transform 1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_85
timestamp 1
transform 1 0 8924 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_89
timestamp 1
transform 1 0 9292 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_93
timestamp 1636968456
transform 1 0 9660 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_132
timestamp 1
transform 1 0 13248 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_138
timestamp 1
transform 1 0 13800 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1636968456
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_153
timestamp 1
transform 1 0 15180 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_10_164
timestamp 1
transform 1 0 16192 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_220
timestamp 1
transform 1 0 21344 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_231
timestamp 1
transform 1 0 22356 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_261
timestamp 1636968456
transform 1 0 25116 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_273
timestamp 1636968456
transform 1 0 26220 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_285
timestamp 1
transform 1 0 27324 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1636968456
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1636968456
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1636968456
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_39
timestamp 1
transform 1 0 4692 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_43
timestamp 1
transform 1 0 5060 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_47
timestamp 1
transform 1 0 5428 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_51
timestamp 1
transform 1 0 5796 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_64
timestamp 1
transform 1 0 6992 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_72
timestamp 1
transform 1 0 7728 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_80
timestamp 1
transform 1 0 8464 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_88
timestamp 1
transform 1 0 9200 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_97
timestamp 1636968456
transform 1 0 10028 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_109
timestamp 1
transform 1 0 11132 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_113
timestamp 1
transform 1 0 11500 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_117
timestamp 1
transform 1 0 11868 0 -1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_11_128
timestamp 1636968456
transform 1 0 12880 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_140
timestamp 1
transform 1 0 13984 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_149
timestamp 1636968456
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_169
timestamp 1
transform 1 0 16652 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_177
timestamp 1636968456
transform 1 0 17388 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_189
timestamp 1
transform 1 0 18492 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_193
timestamp 1
transform 1 0 18860 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_197
timestamp 1
transform 1 0 19228 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_210
timestamp 1636968456
transform 1 0 20424 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_222
timestamp 1
transform 1 0 21528 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_225
timestamp 1
transform 1 0 21804 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_233
timestamp 1
transform 1 0 22540 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_265
timestamp 1636968456
transform 1 0 25484 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_277
timestamp 1
transform 1 0 26588 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_281
timestamp 1
transform 1 0 26956 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_289
timestamp 1
transform 1 0 27692 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1636968456
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1636968456
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1636968456
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_48
timestamp 1
transform 1 0 5520 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_57
timestamp 1636968456
transform 1 0 6348 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_69
timestamp 1
transform 1 0 7452 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_75
timestamp 1
transform 1 0 8004 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_79
timestamp 1
transform 1 0 8372 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_85
timestamp 1
transform 1 0 8924 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_91
timestamp 1
transform 1 0 9476 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1636968456
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_109
timestamp 1
transform 1 0 11132 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_12_126
timestamp 1
transform 1 0 12696 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1636968456
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1636968456
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_165
timestamp 1
transform 1 0 16284 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_178
timestamp 1636968456
transform 1 0 17480 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_190
timestamp 1
transform 1 0 18584 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1636968456
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_209
timestamp 1636968456
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_221
timestamp 1636968456
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_233
timestamp 1
transform 1 0 22540 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_264
timestamp 1636968456
transform 1 0 25392 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_276
timestamp 1636968456
transform 1 0 26496 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_288
timestamp 1
transform 1 0 27600 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1636968456
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1636968456
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1636968456
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1636968456
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1636968456
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1636968456
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_81
timestamp 1
transform 1 0 8556 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_88
timestamp 1636968456
transform 1 0 9200 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_100
timestamp 1636968456
transform 1 0 10304 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_113
timestamp 1
transform 1 0 11500 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_117
timestamp 1
transform 1 0 11868 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_137
timestamp 1636968456
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_149
timestamp 1636968456
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1636968456
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_181
timestamp 1
transform 1 0 17756 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_190
timestamp 1
transform 1 0 18584 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_195
timestamp 1636968456
transform 1 0 19044 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_207
timestamp 1
transform 1 0 20148 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_220
timestamp 1
transform 1 0 21344 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_234
timestamp 1636968456
transform 1 0 22632 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_246
timestamp 1
transform 1 0 23736 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_255
timestamp 1636968456
transform 1 0 24564 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_267
timestamp 1636968456
transform 1 0 25668 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_281
timestamp 1
transform 1 0 26956 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_289
timestamp 1
transform 1 0 27692 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1636968456
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_15
timestamp 1
transform 1 0 2484 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_23
timestamp 1
transform 1 0 3220 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_39
timestamp 1636968456
transform 1 0 4692 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_51
timestamp 1636968456
transform 1 0 5796 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_63
timestamp 1
transform 1 0 6900 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1636968456
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_109
timestamp 1
transform 1 0 11132 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_113
timestamp 1
transform 1 0 11500 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_149
timestamp 1636968456
transform 1 0 14812 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_161
timestamp 1
transform 1 0 15916 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_174
timestamp 1636968456
transform 1 0 17112 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_186
timestamp 1
transform 1 0 18216 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_194
timestamp 1
transform 1 0 18952 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_205
timestamp 1
transform 1 0 19964 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_231
timestamp 1636968456
transform 1 0 22356 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_243
timestamp 1
transform 1 0 23460 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_256
timestamp 1
transform 1 0 24656 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_280
timestamp 1
transform 1 0 26864 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_288
timestamp 1
transform 1 0 27600 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_3
timestamp 1
transform 1 0 1380 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_13
timestamp 1
transform 1 0 2300 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_25
timestamp 1636968456
transform 1 0 3404 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_37
timestamp 1636968456
transform 1 0 4508 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_49
timestamp 1
transform 1 0 5612 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_64
timestamp 1
transform 1 0 6992 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_73
timestamp 1
transform 1 0 7820 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_84
timestamp 1
transform 1 0 8832 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_99
timestamp 1636968456
transform 1 0 10212 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_123
timestamp 1
transform 1 0 12420 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_134
timestamp 1
transform 1 0 13432 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_148
timestamp 1
transform 1 0 14720 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_157
timestamp 1
transform 1 0 15548 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_161
timestamp 1
transform 1 0 15916 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_186
timestamp 1636968456
transform 1 0 18216 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_198
timestamp 1
transform 1 0 19320 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_206
timestamp 1
transform 1 0 20056 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_225
timestamp 1636968456
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_237
timestamp 1
transform 1 0 22908 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_245
timestamp 1
transform 1 0 23644 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_262
timestamp 1636968456
transform 1 0 25208 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_274
timestamp 1
transform 1 0 26312 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_15_281
timestamp 1
transform 1 0 26956 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_289
timestamp 1
transform 1 0 27692 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1636968456
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_15
timestamp 1
transform 1 0 2484 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_19
timestamp 1
transform 1 0 2852 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_23
timestamp 1
transform 1 0 3220 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_36
timestamp 1
transform 1 0 4416 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_50
timestamp 1636968456
transform 1 0 5704 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_62
timestamp 1
transform 1 0 6808 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_72
timestamp 1636968456
transform 1 0 7728 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_85
timestamp 1
transform 1 0 8924 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_96
timestamp 1
transform 1 0 9936 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_107
timestamp 1
transform 1 0 10948 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_115
timestamp 1
transform 1 0 11684 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_124
timestamp 1
transform 1 0 12512 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_138
timestamp 1
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1636968456
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_153
timestamp 1
transform 1 0 15180 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_186
timestamp 1
transform 1 0 18216 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_192
timestamp 1
transform 1 0 18768 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_204
timestamp 1
transform 1 0 19872 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_212
timestamp 1
transform 1 0 20608 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_224
timestamp 1636968456
transform 1 0 21712 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_236
timestamp 1
transform 1 0 22816 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_273
timestamp 1636968456
transform 1 0 26220 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_285
timestamp 1
transform 1 0 27324 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_17_9
timestamp 1636968456
transform 1 0 1932 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_21
timestamp 1
transform 1 0 3036 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_27
timestamp 1
transform 1 0 3588 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_48
timestamp 1
transform 1 0 5520 0 -1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1636968456
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_69
timestamp 1
transform 1 0 7452 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_77
timestamp 1
transform 1 0 8188 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_88
timestamp 1
transform 1 0 9200 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_96
timestamp 1
transform 1 0 9936 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_104
timestamp 1
transform 1 0 10672 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_113
timestamp 1
transform 1 0 11500 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_121
timestamp 1
transform 1 0 12236 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_137
timestamp 1
transform 1 0 13708 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_145
timestamp 1
transform 1 0 14444 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_150
timestamp 1
transform 1 0 14904 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_169
timestamp 1
transform 1 0 16652 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_197
timestamp 1
transform 1 0 19228 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_212
timestamp 1636968456
transform 1 0 20608 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_225
timestamp 1636968456
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_237
timestamp 1
transform 1 0 22908 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_17_256
timestamp 1
transform 1 0 24656 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_262
timestamp 1
transform 1 0 25208 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_269
timestamp 1
transform 1 0 25852 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_277
timestamp 1
transform 1 0 26588 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_281
timestamp 1
transform 1 0 26956 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_289
timestamp 1
transform 1 0 27692 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_3
timestamp 1
transform 1 0 1380 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_20
timestamp 1
transform 1 0 2944 0 1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1636968456
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1636968456
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_53
timestamp 1
transform 1 0 5980 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_70
timestamp 1636968456
transform 1 0 7544 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_82
timestamp 1
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1636968456
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1636968456
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1636968456
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_121
timestamp 1
transform 1 0 12236 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_129
timestamp 1
transform 1 0 12972 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_137
timestamp 1
transform 1 0 13708 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1636968456
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_153
timestamp 1
transform 1 0 15180 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_172
timestamp 1
transform 1 0 16928 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_193
timestamp 1
transform 1 0 18860 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_205
timestamp 1
transform 1 0 19964 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_228
timestamp 1636968456
transform 1 0 22080 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_240
timestamp 1636968456
transform 1 0 23184 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_253
timestamp 1636968456
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_265
timestamp 1636968456
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_277
timestamp 1636968456
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_289
timestamp 1
transform 1 0 27692 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_3
timestamp 1
transform 1 0 1380 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_11
timestamp 1
transform 1 0 2116 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1636968456
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1636968456
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_39
timestamp 1
transform 1 0 4692 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_60
timestamp 1
transform 1 0 6624 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_19_82
timestamp 1
transform 1 0 8648 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_98
timestamp 1636968456
transform 1 0 10120 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_110
timestamp 1
transform 1 0 11224 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1636968456
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_125
timestamp 1
transform 1 0 12604 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_134
timestamp 1636968456
transform 1 0 13432 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_146
timestamp 1
transform 1 0 14536 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_160
timestamp 1
transform 1 0 15824 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_166
timestamp 1
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_169
timestamp 1
transform 1 0 16652 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_178
timestamp 1636968456
transform 1 0 17480 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_193
timestamp 1
transform 1 0 18860 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_201
timestamp 1
transform 1 0 19596 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_219
timestamp 1
transform 1 0 21252 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_235
timestamp 1
transform 1 0 22724 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_252
timestamp 1636968456
transform 1 0 24288 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_264
timestamp 1636968456
transform 1 0 25392 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_276
timestamp 1
transform 1 0 26496 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_281
timestamp 1
transform 1 0 26956 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_289
timestamp 1
transform 1 0 27692 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1636968456
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_15
timestamp 1
transform 1 0 2484 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_29
timestamp 1
transform 1 0 3772 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_46
timestamp 1636968456
transform 1 0 5336 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_58
timestamp 1
transform 1 0 6440 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_62
timestamp 1
transform 1 0 6808 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_67
timestamp 1
transform 1 0 7268 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_75
timestamp 1
transform 1 0 8004 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_101
timestamp 1636968456
transform 1 0 10396 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_113
timestamp 1
transform 1 0 11500 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_122
timestamp 1
transform 1 0 12328 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_133
timestamp 1
transform 1 0 13340 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_141
timestamp 1
transform 1 0 14076 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_20_170
timestamp 1636968456
transform 1 0 16744 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_182
timestamp 1
transform 1 0 17848 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_192
timestamp 1
transform 1 0 18768 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_197
timestamp 1
transform 1 0 19228 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_232
timestamp 1
transform 1 0 22448 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_241
timestamp 1
transform 1 0 23276 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_249
timestamp 1
transform 1 0 24012 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_260
timestamp 1636968456
transform 1 0 25024 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_272
timestamp 1636968456
transform 1 0 26128 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_284
timestamp 1
transform 1 0 27232 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_290
timestamp 1
transform 1 0 27784 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_9
timestamp 1
transform 1 0 1932 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_17
timestamp 1
transform 1 0 2668 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_31
timestamp 1
transform 1 0 3956 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_36
timestamp 1636968456
transform 1 0 4416 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_48
timestamp 1
transform 1 0 5520 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_57
timestamp 1
transform 1 0 6348 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_21_71
timestamp 1
transform 1 0 7636 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_79
timestamp 1
transform 1 0 8372 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_94
timestamp 1636968456
transform 1 0 9752 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_106
timestamp 1
transform 1 0 10856 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_143
timestamp 1
transform 1 0 14260 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_164
timestamp 1
transform 1 0 16192 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_169
timestamp 1
transform 1 0 16652 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_178
timestamp 1
transform 1 0 17480 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_225
timestamp 1
transform 1 0 21804 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_268
timestamp 1636968456
transform 1 0 25760 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_281
timestamp 1
transform 1 0 26956 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_289
timestamp 1
transform 1 0 27692 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1636968456
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_36
timestamp 1
transform 1 0 4416 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_22_68
timestamp 1636968456
transform 1 0 7360 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_80
timestamp 1
transform 1 0 8464 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1636968456
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_97
timestamp 1
transform 1 0 10028 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_105
timestamp 1
transform 1 0 10764 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_141
timestamp 1
transform 1 0 14076 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_164
timestamp 1
transform 1 0 16192 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_168
timestamp 1
transform 1 0 16560 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_176
timestamp 1636968456
transform 1 0 17296 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_188
timestamp 1
transform 1 0 18400 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_22_197
timestamp 1
transform 1 0 19228 0 1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_22_211
timestamp 1636968456
transform 1 0 20516 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_223
timestamp 1636968456
transform 1 0 21620 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_235
timestamp 1
transform 1 0 22724 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_239
timestamp 1
transform 1 0 23092 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_246
timestamp 1
transform 1 0 23736 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_22_266
timestamp 1636968456
transform 1 0 25576 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_278
timestamp 1
transform 1 0 26680 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_286
timestamp 1
transform 1 0 27416 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1636968456
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_15
timestamp 1
transform 1 0 2484 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_21
timestamp 1
transform 1 0 3036 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_26
timestamp 1636968456
transform 1 0 3496 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_38
timestamp 1
transform 1 0 4600 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_46
timestamp 1
transform 1 0 5336 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_53
timestamp 1
transform 1 0 5980 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1636968456
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_69
timestamp 1
transform 1 0 7452 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_73
timestamp 1
transform 1 0 7820 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_96
timestamp 1636968456
transform 1 0 9936 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_108
timestamp 1
transform 1 0 11040 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_132
timestamp 1636968456
transform 1 0 13248 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_144
timestamp 1
transform 1 0 14352 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_23_159
timestamp 1
transform 1 0 15732 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_169
timestamp 1636968456
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_181
timestamp 1
transform 1 0 17756 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_187
timestamp 1
transform 1 0 18308 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_194
timestamp 1636968456
transform 1 0 18952 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_206
timestamp 1
transform 1 0 20056 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_221
timestamp 1
transform 1 0 21436 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_225
timestamp 1636968456
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_237
timestamp 1636968456
transform 1 0 22908 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_249
timestamp 1
transform 1 0 24012 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_253
timestamp 1636968456
transform 1 0 24380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_265
timestamp 1636968456
transform 1 0 25484 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_277
timestamp 1
transform 1 0 26588 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_23_281
timestamp 1
transform 1 0 26956 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_289
timestamp 1
transform 1 0 27692 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_9
timestamp 1
transform 1 0 1932 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_26
timestamp 1
transform 1 0 3496 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_29
timestamp 1
transform 1 0 3772 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_33
timestamp 1
transform 1 0 4140 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_44
timestamp 1636968456
transform 1 0 5152 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_56
timestamp 1636968456
transform 1 0 6256 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_68
timestamp 1
transform 1 0 7360 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_77
timestamp 1
transform 1 0 8188 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_85
timestamp 1
transform 1 0 8924 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_24_110
timestamp 1636968456
transform 1 0 11224 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_122
timestamp 1636968456
transform 1 0 12328 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_134
timestamp 1
transform 1 0 13432 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1636968456
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_153
timestamp 1636968456
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_165
timestamp 1636968456
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_177
timestamp 1636968456
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_189
timestamp 1
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_204
timestamp 1
transform 1 0 19872 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_208
timestamp 1
transform 1 0 20240 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_227
timestamp 1
transform 1 0 21988 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_235
timestamp 1
transform 1 0 22724 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_241
timestamp 1
transform 1 0 23276 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_262
timestamp 1636968456
transform 1 0 25208 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_274
timestamp 1636968456
transform 1 0 26312 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_286
timestamp 1
transform 1 0 27416 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_290
timestamp 1
transform 1 0 27784 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_3
timestamp 1
transform 1 0 1380 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_13
timestamp 1636968456
transform 1 0 2300 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_25
timestamp 1
transform 1 0 3404 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_29
timestamp 1
transform 1 0 3772 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_47
timestamp 1
transform 1 0 5428 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_57
timestamp 1
transform 1 0 6348 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_80
timestamp 1
transform 1 0 8464 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1636968456
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_125
timestamp 1
transform 1 0 12604 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_133
timestamp 1636968456
transform 1 0 13340 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_145
timestamp 1636968456
transform 1 0 14444 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_157
timestamp 1
transform 1 0 15548 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_165
timestamp 1
transform 1 0 16284 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_169
timestamp 1
transform 1 0 16652 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_177
timestamp 1
transform 1 0 17388 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_190
timestamp 1
transform 1 0 18584 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_218
timestamp 1
transform 1 0 21160 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_222
timestamp 1
transform 1 0 21528 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_225
timestamp 1
transform 1 0 21804 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_231
timestamp 1
transform 1 0 22356 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_251
timestamp 1
transform 1 0 24196 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_259
timestamp 1
transform 1 0 24932 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_268
timestamp 1636968456
transform 1 0 25760 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_281
timestamp 1
transform 1 0 26956 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_289
timestamp 1
transform 1 0 27692 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_3
timestamp 1
transform 1 0 1380 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_16
timestamp 1
transform 1 0 2576 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_26
timestamp 1
transform 1 0 3496 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_42
timestamp 1
transform 1 0 4968 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_68
timestamp 1
transform 1 0 7360 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_26_76
timestamp 1
transform 1 0 8096 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_85
timestamp 1
transform 1 0 8924 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_90
timestamp 1636968456
transform 1 0 9384 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_102
timestamp 1636968456
transform 1 0 10488 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_114
timestamp 1
transform 1 0 11592 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_118
timestamp 1
transform 1 0 11960 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_135
timestamp 1
transform 1 0 13524 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1636968456
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_153
timestamp 1636968456
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_165
timestamp 1
transform 1 0 16284 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_173
timestamp 1
transform 1 0 17020 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_194
timestamp 1
transform 1 0 18952 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_197
timestamp 1636968456
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_209
timestamp 1
transform 1 0 20332 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_223
timestamp 1
transform 1 0 21620 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_227
timestamp 1
transform 1 0 21988 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_231
timestamp 1
transform 1 0 22356 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_239
timestamp 1
transform 1 0 23092 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_244
timestamp 1
transform 1 0 23552 0 1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_26_279
timestamp 1636968456
transform 1 0 26772 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_25
timestamp 1
transform 1 0 3404 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_32
timestamp 1636968456
transform 1 0 4048 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_44
timestamp 1636968456
transform 1 0 5152 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_107
timestamp 1
transform 1 0 10948 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_113
timestamp 1
transform 1 0 11500 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_142
timestamp 1
transform 1 0 14168 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_178
timestamp 1
transform 1 0 17480 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_228
timestamp 1636968456
transform 1 0 22080 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_259
timestamp 1636968456
transform 1 0 24932 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_271
timestamp 1
transform 1 0 26036 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_281
timestamp 1
transform 1 0 26956 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_289
timestamp 1
transform 1 0 27692 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_3
timestamp 1
transform 1 0 1380 0 1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1636968456
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1636968456
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1636968456
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_53
timestamp 1
transform 1 0 5980 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_59
timestamp 1
transform 1 0 6532 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_82
timestamp 1
transform 1 0 8648 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_111
timestamp 1636968456
transform 1 0 11316 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_137
timestamp 1
transform 1 0 13708 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_28_141
timestamp 1
transform 1 0 14076 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_28_179
timestamp 1
transform 1 0 17572 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_194
timestamp 1
transform 1 0 18952 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_197
timestamp 1
transform 1 0 19228 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_205
timestamp 1
transform 1 0 19964 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_222
timestamp 1
transform 1 0 21528 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_230
timestamp 1
transform 1 0 22264 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_241
timestamp 1
transform 1 0 23276 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_276
timestamp 1636968456
transform 1 0 26496 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_288
timestamp 1
transform 1 0 27600 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1636968456
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_15
timestamp 1
transform 1 0 2484 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_29_34
timestamp 1
transform 1 0 4232 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_52
timestamp 1
transform 1 0 5888 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_60
timestamp 1
transform 1 0 6624 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_74
timestamp 1636968456
transform 1 0 7912 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_93
timestamp 1
transform 1 0 9660 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_108
timestamp 1
transform 1 0 11040 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 1636968456
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_140
timestamp 1
transform 1 0 13984 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_148
timestamp 1
transform 1 0 14720 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_169
timestamp 1
transform 1 0 16652 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_177
timestamp 1
transform 1 0 17388 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_184
timestamp 1636968456
transform 1 0 18032 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_196
timestamp 1636968456
transform 1 0 19136 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_208
timestamp 1636968456
transform 1 0 20240 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_220
timestamp 1
transform 1 0 21344 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_225
timestamp 1
transform 1 0 21804 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_233
timestamp 1
transform 1 0 22540 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_256
timestamp 1636968456
transform 1 0 24656 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_268
timestamp 1636968456
transform 1 0 25760 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_281
timestamp 1
transform 1 0 26956 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_289
timestamp 1
transform 1 0 27692 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1636968456
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_15
timestamp 1
transform 1 0 2484 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_23
timestamp 1
transform 1 0 3220 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_29
timestamp 1
transform 1 0 3772 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_33
timestamp 1
transform 1 0 4140 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_73
timestamp 1
transform 1 0 7820 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_30_81
timestamp 1
transform 1 0 8556 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_88
timestamp 1
transform 1 0 9200 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_99
timestamp 1636968456
transform 1 0 10212 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_111
timestamp 1636968456
transform 1 0 11316 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_123
timestamp 1
transform 1 0 12420 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_127
timestamp 1
transform 1 0 12788 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_141
timestamp 1
transform 1 0 14076 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_30_156
timestamp 1
transform 1 0 15456 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_30_162
timestamp 1636968456
transform 1 0 16008 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_174
timestamp 1
transform 1 0 17112 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_197
timestamp 1636968456
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_209
timestamp 1
transform 1 0 20332 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_215
timestamp 1
transform 1 0 20884 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_236
timestamp 1636968456
transform 1 0 22816 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_248
timestamp 1
transform 1 0 23920 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_253
timestamp 1636968456
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_265
timestamp 1
transform 1 0 25484 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_22
timestamp 1
transform 1 0 3128 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_47
timestamp 1
transform 1 0 5428 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1636968456
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_69
timestamp 1
transform 1 0 7452 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_87
timestamp 1636968456
transform 1 0 9108 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_99
timestamp 1636968456
transform 1 0 10212 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_113
timestamp 1636968456
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_125
timestamp 1
transform 1 0 12604 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_31_138
timestamp 1636968456
transform 1 0 13800 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_150
timestamp 1636968456
transform 1 0 14904 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_162
timestamp 1
transform 1 0 16008 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_31_169
timestamp 1636968456
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_181
timestamp 1
transform 1 0 17756 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_187
timestamp 1
transform 1 0 18308 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_31_194
timestamp 1
transform 1 0 18952 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_203
timestamp 1636968456
transform 1 0 19780 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_215
timestamp 1
transform 1 0 20884 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_225
timestamp 1
transform 1 0 21804 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_231
timestamp 1
transform 1 0 22356 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_245
timestamp 1636968456
transform 1 0 23644 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_257
timestamp 1636968456
transform 1 0 24748 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_269
timestamp 1
transform 1 0 25852 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_277
timestamp 1
transform 1 0 26588 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_31_281
timestamp 1
transform 1 0 26956 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_9
timestamp 1
transform 1 0 1932 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_26
timestamp 1
transform 1 0 3496 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_29
timestamp 1
transform 1 0 3772 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_33
timestamp 1
transform 1 0 4140 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_37
timestamp 1636968456
transform 1 0 4508 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_49
timestamp 1636968456
transform 1 0 5612 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_61
timestamp 1
transform 1 0 6716 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_67
timestamp 1
transform 1 0 7268 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_75
timestamp 1
transform 1 0 8004 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_98
timestamp 1
transform 1 0 10120 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_141
timestamp 1
transform 1 0 14076 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_147
timestamp 1
transform 1 0 14628 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_151
timestamp 1
transform 1 0 14996 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_157
timestamp 1
transform 1 0 15548 0 1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_32_169
timestamp 1636968456
transform 1 0 16652 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_181
timestamp 1
transform 1 0 17756 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_197
timestamp 1
transform 1 0 19228 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_32_212
timestamp 1
transform 1 0 20608 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_220
timestamp 1
transform 1 0 21344 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_250
timestamp 1
transform 1 0 24104 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_253
timestamp 1636968456
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_265
timestamp 1
transform 1 0 25484 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_286
timestamp 1
transform 1 0 27416 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_290
timestamp 1
transform 1 0 27784 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_33_3
timestamp 1
transform 1 0 1380 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_19
timestamp 1636968456
transform 1 0 2852 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_31
timestamp 1
transform 1 0 3956 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_39
timestamp 1
transform 1 0 4692 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_57
timestamp 1
transform 1 0 6348 0 -1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_33_74
timestamp 1636968456
transform 1 0 7912 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_86
timestamp 1636968456
transform 1 0 9016 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_98
timestamp 1636968456
transform 1 0 10120 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_110
timestamp 1
transform 1 0 11224 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_128
timestamp 1
transform 1 0 12880 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_143
timestamp 1
transform 1 0 14260 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_33_221
timestamp 1
transform 1 0 21436 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_253
timestamp 1636968456
transform 1 0 24380 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_265
timestamp 1
transform 1 0 25484 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_278
timestamp 1
transform 1 0 26680 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_281
timestamp 1
transform 1 0 26956 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_289
timestamp 1
transform 1 0 27692 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_15
timestamp 1636968456
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_32
timestamp 1
transform 1 0 4048 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_43
timestamp 1
transform 1 0 5060 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_53
timestamp 1
transform 1 0 5980 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_34_66
timestamp 1636968456
transform 1 0 7176 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_78
timestamp 1
transform 1 0 8280 0 1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 1636968456
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_97
timestamp 1
transform 1 0 10028 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_34_147
timestamp 1
transform 1 0 14628 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_162
timestamp 1
transform 1 0 16008 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_173
timestamp 1
transform 1 0 17020 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_182
timestamp 1
transform 1 0 17848 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_34_194
timestamp 1
transform 1 0 18952 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_245
timestamp 1
transform 1 0 23644 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 1
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_253
timestamp 1
transform 1 0 24380 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_257
timestamp 1
transform 1 0 24748 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_283
timestamp 1
transform 1 0 27140 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_3
timestamp 1
transform 1 0 1380 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_19
timestamp 1
transform 1 0 2852 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_23
timestamp 1
transform 1 0 3220 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_50
timestamp 1
transform 1 0 5704 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_35_57
timestamp 1
transform 1 0 6348 0 -1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_35_78
timestamp 1636968456
transform 1 0 8280 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_90
timestamp 1636968456
transform 1 0 9384 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_102
timestamp 1
transform 1 0 10488 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_110
timestamp 1
transform 1 0 11224 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_113
timestamp 1636968456
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_146
timestamp 1
transform 1 0 14536 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_155
timestamp 1
transform 1 0 15364 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_161
timestamp 1
transform 1 0 15916 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_169
timestamp 1
transform 1 0 16652 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_173
timestamp 1
transform 1 0 17020 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_196
timestamp 1
transform 1 0 19136 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_200
timestamp 1
transform 1 0 19504 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_205
timestamp 1
transform 1 0 19964 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_212
timestamp 1636968456
transform 1 0 20608 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_225
timestamp 1
transform 1 0 21804 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_233
timestamp 1
transform 1 0 22540 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_241
timestamp 1636968456
transform 1 0 23276 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_253
timestamp 1
transform 1 0 24380 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_35_277
timestamp 1
transform 1 0 26588 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_35_285
timestamp 1
transform 1 0 27324 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_6
timestamp 1
transform 1 0 1656 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_24
timestamp 1
transform 1 0 3312 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_39
timestamp 1636968456
transform 1 0 4692 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_51
timestamp 1636968456
transform 1 0 5796 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_63
timestamp 1
transform 1 0 6900 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_70
timestamp 1636968456
transform 1 0 7544 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_82
timestamp 1
transform 1 0 8648 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_85
timestamp 1
transform 1 0 8924 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_36_104
timestamp 1636968456
transform 1 0 10672 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_116
timestamp 1636968456
transform 1 0 11776 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_128
timestamp 1
transform 1 0 12880 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_132
timestamp 1
transform 1 0 13248 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_136
timestamp 1
transform 1 0 13616 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_141
timestamp 1
transform 1 0 14076 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_36_157
timestamp 1
transform 1 0 15548 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_163
timestamp 1
transform 1 0 16100 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_179
timestamp 1636968456
transform 1 0 17572 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_191
timestamp 1
transform 1 0 18676 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_197
timestamp 1636968456
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_209
timestamp 1636968456
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_221
timestamp 1636968456
transform 1 0 21436 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_233
timestamp 1636968456
transform 1 0 22540 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_245
timestamp 1
transform 1 0 23644 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_253
timestamp 1
transform 1 0 24380 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_261
timestamp 1
transform 1 0 25116 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_275
timestamp 1636968456
transform 1 0 26404 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_287
timestamp 1
transform 1 0 27508 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_7
timestamp 1
transform 1 0 1748 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_11
timestamp 1
transform 1 0 2116 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_31
timestamp 1636968456
transform 1 0 3956 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_43
timestamp 1
transform 1 0 5060 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_37_53
timestamp 1
transform 1 0 5980 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_37_57
timestamp 1
transform 1 0 6348 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_61
timestamp 1
transform 1 0 6716 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_69
timestamp 1
transform 1 0 7452 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_77
timestamp 1
transform 1 0 8188 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_81
timestamp 1
transform 1 0 8556 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_87
timestamp 1
transform 1 0 9108 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_101
timestamp 1
transform 1 0 10396 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_109
timestamp 1
transform 1 0 11132 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_37_113
timestamp 1636968456
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_125
timestamp 1
transform 1 0 12604 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_137
timestamp 1
transform 1 0 13708 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_146
timestamp 1636968456
transform 1 0 14536 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_158
timestamp 1
transform 1 0 15640 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_166
timestamp 1
transform 1 0 16376 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_169
timestamp 1
transform 1 0 16652 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_179
timestamp 1636968456
transform 1 0 17572 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_191
timestamp 1
transform 1 0 18676 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_195
timestamp 1
transform 1 0 19044 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_203
timestamp 1
transform 1 0 19780 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_211
timestamp 1
transform 1 0 20516 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_222
timestamp 1
transform 1 0 21528 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_225
timestamp 1636968456
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_237
timestamp 1636968456
transform 1 0 22908 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_249
timestamp 1636968456
transform 1 0 24012 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_261
timestamp 1
transform 1 0 25116 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_268
timestamp 1
transform 1 0 25760 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_272
timestamp 1
transform 1 0 26128 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_277
timestamp 1
transform 1 0 26588 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_37_286
timestamp 1
transform 1 0 27416 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1636968456
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1636968456
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_29
timestamp 1
transform 1 0 3772 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_33
timestamp 1
transform 1 0 4140 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_37
timestamp 1
transform 1 0 4508 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_52
timestamp 1
transform 1 0 5888 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_78
timestamp 1
transform 1 0 8280 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_38_85
timestamp 1
transform 1 0 8924 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_108
timestamp 1636968456
transform 1 0 11040 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_120
timestamp 1
transform 1 0 12144 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_135
timestamp 1
transform 1 0 13524 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_141
timestamp 1636968456
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_153
timestamp 1636968456
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_165
timestamp 1636968456
transform 1 0 16284 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_177
timestamp 1636968456
transform 1 0 17388 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_197
timestamp 1
transform 1 0 19228 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_213
timestamp 1636968456
transform 1 0 20700 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_225
timestamp 1
transform 1 0 21804 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_231
timestamp 1
transform 1 0 22356 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_242
timestamp 1
transform 1 0 23368 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_248
timestamp 1
transform 1 0 23920 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_273
timestamp 1
transform 1 0 26220 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_281
timestamp 1
transform 1 0 26956 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_289
timestamp 1
transform 1 0 27692 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_28
timestamp 1
transform 1 0 3680 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_39_50
timestamp 1
transform 1 0 5704 0 -1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1636968456
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_69
timestamp 1636968456
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_39_81
timestamp 1
transform 1 0 8556 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_87
timestamp 1
transform 1 0 9108 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_96
timestamp 1636968456
transform 1 0 9936 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_108
timestamp 1
transform 1 0 11040 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_113
timestamp 1
transform 1 0 11500 0 -1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_39_134
timestamp 1636968456
transform 1 0 13432 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_146
timestamp 1636968456
transform 1 0 14536 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_158
timestamp 1
transform 1 0 15640 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_39_162
timestamp 1
transform 1 0 16008 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_186
timestamp 1
transform 1 0 18216 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_196
timestamp 1
transform 1 0 19136 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_203
timestamp 1636968456
transform 1 0 19780 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_215
timestamp 1
transform 1 0 20884 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_248
timestamp 1
transform 1 0 23920 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_256
timestamp 1
transform 1 0 24656 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_269
timestamp 1
transform 1 0 25852 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_277
timestamp 1
transform 1 0 26588 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_39_281
timestamp 1
transform 1 0 26956 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_40_22
timestamp 1
transform 1 0 3128 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_40_48
timestamp 1636968456
transform 1 0 5520 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_60
timestamp 1
transform 1 0 6624 0 1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_40_71
timestamp 1636968456
transform 1 0 7636 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_103
timestamp 1636968456
transform 1 0 10580 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_115
timestamp 1
transform 1 0 11684 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_138
timestamp 1
transform 1 0 13800 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_146
timestamp 1
transform 1 0 14536 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_40_189
timestamp 1
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_218
timestamp 1
transform 1 0 21160 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_257
timestamp 1
transform 1 0 24748 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_3
timestamp 1636968456
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_15
timestamp 1636968456
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_27
timestamp 1
transform 1 0 3588 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_31
timestamp 1
transform 1 0 3956 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_39
timestamp 1636968456
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1636968456
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_69
timestamp 1
transform 1 0 7452 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_73
timestamp 1
transform 1 0 7820 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_88
timestamp 1
transform 1 0 9200 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_94
timestamp 1
transform 1 0 9752 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_108
timestamp 1
transform 1 0 11040 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_113
timestamp 1
transform 1 0 11500 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_132
timestamp 1636968456
transform 1 0 13248 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_144
timestamp 1
transform 1 0 14352 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_150
timestamp 1
transform 1 0 14904 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_161
timestamp 1
transform 1 0 15916 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_180
timestamp 1636968456
transform 1 0 17664 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_192
timestamp 1636968456
transform 1 0 18768 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_204
timestamp 1636968456
transform 1 0 19872 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_216
timestamp 1
transform 1 0 20976 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_225
timestamp 1
transform 1 0 21804 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_250
timestamp 1636968456
transform 1 0 24104 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_41_284
timestamp 1
transform 1 0 27232 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_42_3
timestamp 1
transform 1 0 1380 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_11
timestamp 1
transform 1 0 2116 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_26
timestamp 1
transform 1 0 3496 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1636968456
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1636968456
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_53
timestamp 1
transform 1 0 5980 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_42_69
timestamp 1
transform 1 0 7452 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_73
timestamp 1
transform 1 0 7820 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_42_78
timestamp 1
transform 1 0 8280 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_85
timestamp 1
transform 1 0 8924 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_92
timestamp 1
transform 1 0 9568 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_96
timestamp 1
transform 1 0 9936 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_102
timestamp 1636968456
transform 1 0 10488 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_114
timestamp 1
transform 1 0 11592 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_42_129
timestamp 1
transform 1 0 12972 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_137
timestamp 1
transform 1 0 13708 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_42_141
timestamp 1
transform 1 0 14076 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_149
timestamp 1
transform 1 0 14812 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_42_166
timestamp 1636968456
transform 1 0 16376 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_178
timestamp 1636968456
transform 1 0 17480 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_190
timestamp 1
transform 1 0 18584 0 1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_42_197
timestamp 1636968456
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_209
timestamp 1
transform 1 0 20332 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_219
timestamp 1636968456
transform 1 0 21252 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_231
timestamp 1
transform 1 0 22356 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_245
timestamp 1
transform 1 0 23644 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_253
timestamp 1636968456
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_265
timestamp 1
transform 1 0 25484 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_42_284
timestamp 1
transform 1 0 27232 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1636968456
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_15
timestamp 1
transform 1 0 2484 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_23
timestamp 1636968456
transform 1 0 3220 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_35
timestamp 1636968456
transform 1 0 4324 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_47
timestamp 1
transform 1 0 5428 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1636968456
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_43_69
timestamp 1
transform 1 0 7452 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_43_77
timestamp 1636968456
transform 1 0 8188 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_89
timestamp 1636968456
transform 1 0 9292 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_104
timestamp 1
transform 1 0 10672 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_43_113
timestamp 1
transform 1 0 11500 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_121
timestamp 1
transform 1 0 12236 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_43_127
timestamp 1636968456
transform 1 0 12788 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_139
timestamp 1636968456
transform 1 0 13892 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_151
timestamp 1636968456
transform 1 0 14996 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_163
timestamp 1
transform 1 0 16100 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_169
timestamp 1636968456
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_181
timestamp 1636968456
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_193
timestamp 1636968456
transform 1 0 18860 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_205
timestamp 1636968456
transform 1 0 19964 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_217
timestamp 1
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_225
timestamp 1636968456
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_237
timestamp 1636968456
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_249
timestamp 1636968456
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_261
timestamp 1636968456
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_278
timestamp 1
transform 1 0 26680 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_43_284
timestamp 1
transform 1 0 27232 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_290
timestamp 1
transform 1 0 27784 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_44_3
timestamp 1
transform 1 0 1380 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_23
timestamp 1
transform 1 0 3220 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_32
timestamp 1
transform 1 0 4048 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_40
timestamp 1
transform 1 0 4784 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_44_52
timestamp 1
transform 1 0 5888 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_44_66
timestamp 1
transform 1 0 7176 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_44_72
timestamp 1
transform 1 0 7728 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_91
timestamp 1
transform 1 0 9476 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_44_110
timestamp 1
transform 1 0 11224 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_118
timestamp 1
transform 1 0 11960 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_135
timestamp 1
transform 1 0 13524 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_141
timestamp 1636968456
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_153
timestamp 1636968456
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_165
timestamp 1636968456
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_177
timestamp 1636968456
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_189
timestamp 1
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_197
timestamp 1
transform 1 0 19228 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_211
timestamp 1
transform 1 0 20516 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_218
timestamp 1636968456
transform 1 0 21160 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_230
timestamp 1
transform 1 0 22264 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_234
timestamp 1
transform 1 0 22632 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_240
timestamp 1636968456
transform 1 0 23184 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_253
timestamp 1
transform 1 0 24380 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_257
timestamp 1
transform 1 0 24748 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_44_269
timestamp 1
transform 1 0 25852 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_280
timestamp 1
transform 1 0 26864 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_286
timestamp 1
transform 1 0 27416 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_3
timestamp 1
transform 1 0 1380 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_9
timestamp 1
transform 1 0 1932 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_45_17
timestamp 1
transform 1 0 2668 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_45_36
timestamp 1
transform 1 0 4416 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_57
timestamp 1
transform 1 0 6348 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_71
timestamp 1636968456
transform 1 0 7636 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_90
timestamp 1
transform 1 0 9384 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_100
timestamp 1
transform 1 0 10304 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_127
timestamp 1636968456
transform 1 0 12788 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_139
timestamp 1636968456
transform 1 0 13892 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_151
timestamp 1636968456
transform 1 0 14996 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_163
timestamp 1
transform 1 0 16100 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_169
timestamp 1
transform 1 0 16652 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_175
timestamp 1
transform 1 0 17204 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_45_179
timestamp 1
transform 1 0 17572 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_45_222
timestamp 1
transform 1 0 21528 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_45_235
timestamp 1
transform 1 0 22724 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_241
timestamp 1
transform 1 0 23276 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_249
timestamp 1
transform 1 0 24012 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_261
timestamp 1
transform 1 0 25116 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_45_266
timestamp 1
transform 1 0 25576 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_275
timestamp 1
transform 1 0 26404 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 1
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_281
timestamp 1
transform 1 0 26956 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_289
timestamp 1
transform 1 0 27692 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1636968456
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_15
timestamp 1636968456
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1636968456
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_41
timestamp 1
transform 1 0 4876 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_49
timestamp 1
transform 1 0 5612 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_72
timestamp 1636968456
transform 1 0 7728 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_85
timestamp 1
transform 1 0 8924 0 1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_46_118
timestamp 1636968456
transform 1 0 11960 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_130
timestamp 1
transform 1 0 13064 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_138
timestamp 1
transform 1 0 13800 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_141
timestamp 1636968456
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_153
timestamp 1636968456
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_165
timestamp 1
transform 1 0 16284 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_171
timestamp 1
transform 1 0 16836 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_247
timestamp 1
transform 1 0 23828 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_46_285
timestamp 1
transform 1 0 27324 0 1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_47_3
timestamp 1636968456
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_15
timestamp 1636968456
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_27
timestamp 1636968456
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_39
timestamp 1636968456
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1636968456
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_69
timestamp 1636968456
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_81
timestamp 1636968456
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_93
timestamp 1
transform 1 0 9660 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_99
timestamp 1
transform 1 0 10212 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_113
timestamp 1636968456
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_125
timestamp 1636968456
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_137
timestamp 1636968456
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_149
timestamp 1636968456
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_161
timestamp 1
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_169
timestamp 1636968456
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_181
timestamp 1
transform 1 0 17756 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_192
timestamp 1
transform 1 0 18768 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_47_212
timestamp 1
transform 1 0 20608 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_220
timestamp 1
transform 1 0 21344 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_225
timestamp 1
transform 1 0 21804 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_230
timestamp 1636968456
transform 1 0 22264 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_242
timestamp 1636968456
transform 1 0 23368 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_254
timestamp 1
transform 1 0 24472 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_261
timestamp 1636968456
transform 1 0 25116 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_273
timestamp 1
transform 1 0 26220 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_279
timestamp 1
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_281
timestamp 1
transform 1 0 26956 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1636968456
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_15
timestamp 1636968456
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1636968456
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_41
timestamp 1636968456
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_48_53
timestamp 1
transform 1 0 5980 0 1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_48_57
timestamp 1636968456
transform 1 0 6348 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_69
timestamp 1636968456
transform 1 0 7452 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_48_81
timestamp 1
transform 1 0 8556 0 1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_48_85
timestamp 1636968456
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_97
timestamp 1636968456
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_48_109
timestamp 1
transform 1 0 11132 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_48_113
timestamp 1
transform 1 0 11500 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_48_119
timestamp 1
transform 1 0 12052 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_48_126
timestamp 1
transform 1 0 12696 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_48_133
timestamp 1
transform 1 0 13340 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_48_141
timestamp 1
transform 1 0 14076 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_48_147
timestamp 1
transform 1 0 14628 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_48_154
timestamp 1
transform 1 0 15272 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_48_161
timestamp 1
transform 1 0 15916 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_48_169
timestamp 1
transform 1 0 16652 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_48_175
timestamp 1
transform 1 0 17204 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_48_182
timestamp 1
transform 1 0 17848 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_48_189
timestamp 1
transform 1 0 18492 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_48_197
timestamp 1
transform 1 0 19228 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_48_203
timestamp 1
transform 1 0 19780 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_48_210
timestamp 1
transform 1 0 20424 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_48_217
timestamp 1
transform 1 0 21068 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_48_225
timestamp 1
transform 1 0 21804 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_48_231
timestamp 1
transform 1 0 22356 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_48_238
timestamp 1
transform 1 0 23000 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_48_245
timestamp 1
transform 1 0 23644 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_48_253
timestamp 1
transform 1 0 24380 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_48_259
timestamp 1
transform 1 0 24932 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_48_266
timestamp 1
transform 1 0 25576 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_48_273
timestamp 1
transform 1 0 26220 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_48_281
timestamp 1
transform 1 0 26956 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1
transform 1 0 27600 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1
transform 1 0 27600 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input3
timestamp 1
transform 1 0 9108 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input4
timestamp 1
transform 1 0 1380 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input5
timestamp 1
transform 1 0 1380 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 1
transform 1 0 1380 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input7
timestamp 1
transform 1 0 1380 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input8
timestamp 1
transform 1 0 5888 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  input9
timestamp 1
transform 1 0 1380 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input10
timestamp 1
transform 1 0 1380 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input11
timestamp 1
transform 1 0 1380 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input12
timestamp 1
transform 1 0 1380 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input13
timestamp 1
transform 1 0 1380 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input14
timestamp 1
transform 1 0 1932 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input15
timestamp 1
transform 1 0 1380 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  input16
timestamp 1
transform 1 0 1380 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input17
timestamp 1
transform -1 0 27876 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output18
timestamp 1
transform -1 0 27876 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output19
timestamp 1
transform 1 0 23276 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output20
timestamp 1
transform 1 0 23920 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output21
timestamp 1
transform 1 0 27508 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output22
timestamp 1
transform -1 0 12052 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output23
timestamp 1
transform -1 0 15916 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output24
timestamp 1
transform -1 0 13340 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output25
timestamp 1
transform -1 0 18492 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output26
timestamp 1
transform -1 0 22356 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output27
timestamp 1
transform 1 0 22632 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output28
timestamp 1
transform -1 0 15272 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output29
timestamp 1
transform 1 0 27140 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output30
timestamp 1
transform 1 0 27508 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output31
timestamp 1
transform -1 0 16560 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output32
timestamp 1
transform 1 0 21344 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output33
timestamp 1
transform 1 0 20056 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output34
timestamp 1
transform 1 0 25852 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output35
timestamp 1
transform -1 0 17848 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output36
timestamp 1
transform 1 0 26496 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output37
timestamp 1
transform 1 0 27508 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output38
timestamp 1
transform 1 0 25208 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output39
timestamp 1
transform -1 0 14628 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output40
timestamp 1
transform -1 0 17204 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output41
timestamp 1
transform 1 0 19412 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output42
timestamp 1
transform 1 0 27508 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output43
timestamp 1
transform 1 0 27508 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output44
timestamp 1
transform 1 0 27508 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output45
timestamp 1
transform 1 0 27508 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output46
timestamp 1
transform 1 0 27140 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output47
timestamp 1
transform -1 0 12696 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output48
timestamp 1
transform -1 0 19136 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output49
timestamp 1
transform -1 0 13984 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output50
timestamp 1
transform 1 0 24564 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output51
timestamp 1
transform 1 0 20700 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output52
timestamp 1
transform 1 0 27508 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_49
timestamp 1
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1
transform -1 0 28152 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_50
timestamp 1
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1
transform -1 0 28152 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_51
timestamp 1
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1
transform -1 0 28152 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_52
timestamp 1
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1
transform -1 0 28152 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_53
timestamp 1
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1
transform -1 0 28152 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_54
timestamp 1
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1
transform -1 0 28152 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_55
timestamp 1
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1
transform -1 0 28152 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_56
timestamp 1
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1
transform -1 0 28152 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_57
timestamp 1
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1
transform -1 0 28152 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_58
timestamp 1
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1
transform -1 0 28152 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_59
timestamp 1
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1
transform -1 0 28152 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_60
timestamp 1
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1
transform -1 0 28152 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_61
timestamp 1
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1
transform -1 0 28152 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_62
timestamp 1
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1
transform -1 0 28152 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_63
timestamp 1
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1
transform -1 0 28152 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_64
timestamp 1
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1
transform -1 0 28152 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_65
timestamp 1
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1
transform -1 0 28152 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_66
timestamp 1
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 1
transform -1 0 28152 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_67
timestamp 1
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 1
transform -1 0 28152 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_68
timestamp 1
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 1
transform -1 0 28152 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_69
timestamp 1
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 1
transform -1 0 28152 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_70
timestamp 1
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 1
transform -1 0 28152 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_71
timestamp 1
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 1
transform -1 0 28152 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_72
timestamp 1
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 1
transform -1 0 28152 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_73
timestamp 1
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 1
transform -1 0 28152 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_74
timestamp 1
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 1
transform -1 0 28152 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_75
timestamp 1
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 1
transform -1 0 28152 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_76
timestamp 1
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 1
transform -1 0 28152 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_77
timestamp 1
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 1
transform -1 0 28152 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_78
timestamp 1
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp 1
transform -1 0 28152 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_79
timestamp 1
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp 1
transform -1 0 28152 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_80
timestamp 1
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp 1
transform -1 0 28152 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_81
timestamp 1
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp 1
transform -1 0 28152 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Left_82
timestamp 1
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Right_33
timestamp 1
transform -1 0 28152 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Left_83
timestamp 1
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Right_34
timestamp 1
transform -1 0 28152 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Left_84
timestamp 1
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Right_35
timestamp 1
transform -1 0 28152 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Left_85
timestamp 1
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Right_36
timestamp 1
transform -1 0 28152 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Left_86
timestamp 1
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Right_37
timestamp 1
transform -1 0 28152 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Left_87
timestamp 1
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Right_38
timestamp 1
transform -1 0 28152 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Left_88
timestamp 1
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Right_39
timestamp 1
transform -1 0 28152 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Left_89
timestamp 1
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Right_40
timestamp 1
transform -1 0 28152 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Left_90
timestamp 1
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Right_41
timestamp 1
transform -1 0 28152 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Left_91
timestamp 1
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Right_42
timestamp 1
transform -1 0 28152 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Left_92
timestamp 1
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Right_43
timestamp 1
transform -1 0 28152 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Left_93
timestamp 1
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Right_44
timestamp 1
transform -1 0 28152 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Left_94
timestamp 1
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Right_45
timestamp 1
transform -1 0 28152 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Left_95
timestamp 1
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Right_46
timestamp 1
transform -1 0 28152 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_Left_96
timestamp 1
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_Right_47
timestamp 1
transform -1 0 28152 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_Left_97
timestamp 1
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_Right_48
timestamp 1
transform -1 0 28152 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_98
timestamp 1
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_99
timestamp 1
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_100
timestamp 1
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_101
timestamp 1
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_102
timestamp 1
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_103
timestamp 1
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_104
timestamp 1
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_105
timestamp 1
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_106
timestamp 1
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_107
timestamp 1
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_108
timestamp 1
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_109
timestamp 1
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_110
timestamp 1
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_111
timestamp 1
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_112
timestamp 1
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_113
timestamp 1
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_114
timestamp 1
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_115
timestamp 1
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_116
timestamp 1
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_117
timestamp 1
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_118
timestamp 1
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_119
timestamp 1
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_120
timestamp 1
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_121
timestamp 1
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_122
timestamp 1
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_123
timestamp 1
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_124
timestamp 1
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_125
timestamp 1
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_126
timestamp 1
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_127
timestamp 1
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_128
timestamp 1
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_129
timestamp 1
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_130
timestamp 1
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_131
timestamp 1
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_132
timestamp 1
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_133
timestamp 1
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_134
timestamp 1
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_135
timestamp 1
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_136
timestamp 1
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_137
timestamp 1
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_138
timestamp 1
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_139
timestamp 1
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_140
timestamp 1
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_141
timestamp 1
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_142
timestamp 1
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_143
timestamp 1
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_144
timestamp 1
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_145
timestamp 1
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_146
timestamp 1
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_147
timestamp 1
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_148
timestamp 1
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_149
timestamp 1
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_150
timestamp 1
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_151
timestamp 1
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_152
timestamp 1
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_153
timestamp 1
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_154
timestamp 1
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_155
timestamp 1
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_156
timestamp 1
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_157
timestamp 1
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_158
timestamp 1
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_159
timestamp 1
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_160
timestamp 1
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_161
timestamp 1
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_162
timestamp 1
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_163
timestamp 1
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_164
timestamp 1
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_165
timestamp 1
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_166
timestamp 1
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_167
timestamp 1
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_168
timestamp 1
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_169
timestamp 1
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_170
timestamp 1
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_171
timestamp 1
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_172
timestamp 1
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_173
timestamp 1
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_174
timestamp 1
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_175
timestamp 1
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_176
timestamp 1
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_177
timestamp 1
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_178
timestamp 1
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_179
timestamp 1
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_180
timestamp 1
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_181
timestamp 1
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_182
timestamp 1
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_183
timestamp 1
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_184
timestamp 1
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_185
timestamp 1
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_186
timestamp 1
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_187
timestamp 1
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_188
timestamp 1
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_189
timestamp 1
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_190
timestamp 1
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_191
timestamp 1
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_192
timestamp 1
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_193
timestamp 1
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_194
timestamp 1
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_195
timestamp 1
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_196
timestamp 1
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_197
timestamp 1
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_198
timestamp 1
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_199
timestamp 1
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_200
timestamp 1
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_201
timestamp 1
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_202
timestamp 1
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_203
timestamp 1
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_204
timestamp 1
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_205
timestamp 1
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_206
timestamp 1
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_207
timestamp 1
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_208
timestamp 1
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_209
timestamp 1
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_210
timestamp 1
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_211
timestamp 1
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_212
timestamp 1
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_213
timestamp 1
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_214
timestamp 1
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_215
timestamp 1
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_216
timestamp 1
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_217
timestamp 1
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_218
timestamp 1
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_219
timestamp 1
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_220
timestamp 1
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_221
timestamp 1
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_222
timestamp 1
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_223
timestamp 1
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_224
timestamp 1
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_225
timestamp 1
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_226
timestamp 1
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_227
timestamp 1
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_228
timestamp 1
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_229
timestamp 1
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_230
timestamp 1
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_231
timestamp 1
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_232
timestamp 1
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_233
timestamp 1
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_234
timestamp 1
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_235
timestamp 1
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_236
timestamp 1
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_237
timestamp 1
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_238
timestamp 1
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_239
timestamp 1
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_240
timestamp 1
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_241
timestamp 1
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_242
timestamp 1
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_243
timestamp 1
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_244
timestamp 1
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_245
timestamp 1
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_246
timestamp 1
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_247
timestamp 1
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_248
timestamp 1
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_249
timestamp 1
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_250
timestamp 1
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_251
timestamp 1
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_252
timestamp 1
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_253
timestamp 1
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_254
timestamp 1
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_255
timestamp 1
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_256
timestamp 1
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_257
timestamp 1
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_258
timestamp 1
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_259
timestamp 1
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_260
timestamp 1
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_261
timestamp 1
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_262
timestamp 1
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_263
timestamp 1
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_264
timestamp 1
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_265
timestamp 1
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_266
timestamp 1
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_267
timestamp 1
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_268
timestamp 1
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_269
timestamp 1
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_270
timestamp 1
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_271
timestamp 1
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_272
timestamp 1
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_273
timestamp 1
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_274
timestamp 1
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_275
timestamp 1
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_276
timestamp 1
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_277
timestamp 1
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_278
timestamp 1
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_279
timestamp 1
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_280
timestamp 1
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_281
timestamp 1
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_282
timestamp 1
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_283
timestamp 1
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_284
timestamp 1
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_285
timestamp 1
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_286
timestamp 1
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_287
timestamp 1
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_288
timestamp 1
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_289
timestamp 1
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_290
timestamp 1
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_291
timestamp 1
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_292
timestamp 1
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_293
timestamp 1
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_294
timestamp 1
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_295
timestamp 1
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_296
timestamp 1
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_297
timestamp 1
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_298
timestamp 1
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_299
timestamp 1
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_300
timestamp 1
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_301
timestamp 1
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_302
timestamp 1
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_303
timestamp 1
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_304
timestamp 1
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_305
timestamp 1
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_306
timestamp 1
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_307
timestamp 1
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_308
timestamp 1
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_309
timestamp 1
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_310
timestamp 1
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_311
timestamp 1
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_312
timestamp 1
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_313
timestamp 1
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_314
timestamp 1
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_315
timestamp 1
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_316
timestamp 1
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_317
timestamp 1
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_318
timestamp 1
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_319
timestamp 1
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_320
timestamp 1
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_321
timestamp 1
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_322
timestamp 1
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_323
timestamp 1
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_324
timestamp 1
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_325
timestamp 1
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_326
timestamp 1
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_327
timestamp 1
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_328
timestamp 1
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_329
timestamp 1
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_330
timestamp 1
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_331
timestamp 1
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_332
timestamp 1
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_333
timestamp 1
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_334
timestamp 1
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_335
timestamp 1
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_336
timestamp 1
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_337
timestamp 1
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_338
timestamp 1
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_339
timestamp 1
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_340
timestamp 1
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_341
timestamp 1
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_342
timestamp 1
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_343
timestamp 1
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_344
timestamp 1
transform 1 0 6256 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_345
timestamp 1
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_346
timestamp 1
transform 1 0 11408 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_347
timestamp 1
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_348
timestamp 1
transform 1 0 16560 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_349
timestamp 1
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_350
timestamp 1
transform 1 0 21712 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_351
timestamp 1
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_352
timestamp 1
transform 1 0 26864 0 1 28288
box -38 -48 130 592
<< labels >>
flabel metal4 s 4868 2128 5188 28880 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 4208 2128 4528 28880 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 28532 4768 29332 4888 0 FreeSans 480 0 0 0 clk
port 2 nsew signal input
flabel metal3 s 28532 19048 29332 19168 0 FreeSans 480 0 0 0 done
port 3 nsew signal output
flabel metal3 s 28532 6128 29332 6248 0 FreeSans 480 0 0 0 enable
port 4 nsew signal input
flabel metal3 s 28532 5448 29332 5568 0 FreeSans 480 0 0 0 nrst
port 5 nsew signal input
flabel metal2 s 23202 30676 23258 31476 0 FreeSans 224 90 0 0 out[0]
port 6 nsew signal output
flabel metal2 s 23846 30676 23902 31476 0 FreeSans 224 90 0 0 out[10]
port 7 nsew signal output
flabel metal2 s 28998 30676 29054 31476 0 FreeSans 224 90 0 0 out[11]
port 8 nsew signal output
flabel metal2 s 11610 30676 11666 31476 0 FreeSans 224 90 0 0 out[12]
port 9 nsew signal output
flabel metal2 s 15474 30676 15530 31476 0 FreeSans 224 90 0 0 out[13]
port 10 nsew signal output
flabel metal2 s 12898 30676 12954 31476 0 FreeSans 224 90 0 0 out[14]
port 11 nsew signal output
flabel metal2 s 18050 30676 18106 31476 0 FreeSans 224 90 0 0 out[15]
port 12 nsew signal output
flabel metal2 s 21914 30676 21970 31476 0 FreeSans 224 90 0 0 out[16]
port 13 nsew signal output
flabel metal2 s 22558 30676 22614 31476 0 FreeSans 224 90 0 0 out[17]
port 14 nsew signal output
flabel metal2 s 14830 30676 14886 31476 0 FreeSans 224 90 0 0 out[18]
port 15 nsew signal output
flabel metal2 s 27066 30676 27122 31476 0 FreeSans 224 90 0 0 out[19]
port 16 nsew signal output
flabel metal3 s 28532 24488 29332 24608 0 FreeSans 480 0 0 0 out[1]
port 17 nsew signal output
flabel metal2 s 16118 30676 16174 31476 0 FreeSans 224 90 0 0 out[20]
port 18 nsew signal output
flabel metal2 s 21270 30676 21326 31476 0 FreeSans 224 90 0 0 out[21]
port 19 nsew signal output
flabel metal2 s 19982 30676 20038 31476 0 FreeSans 224 90 0 0 out[22]
port 20 nsew signal output
flabel metal2 s 25778 30676 25834 31476 0 FreeSans 224 90 0 0 out[23]
port 21 nsew signal output
flabel metal2 s 17406 30676 17462 31476 0 FreeSans 224 90 0 0 out[24]
port 22 nsew signal output
flabel metal2 s 26422 30676 26478 31476 0 FreeSans 224 90 0 0 out[25]
port 23 nsew signal output
flabel metal3 s 28532 25848 29332 25968 0 FreeSans 480 0 0 0 out[26]
port 24 nsew signal output
flabel metal2 s 25134 30676 25190 31476 0 FreeSans 224 90 0 0 out[27]
port 25 nsew signal output
flabel metal2 s 14186 30676 14242 31476 0 FreeSans 224 90 0 0 out[28]
port 26 nsew signal output
flabel metal2 s 16762 30676 16818 31476 0 FreeSans 224 90 0 0 out[29]
port 27 nsew signal output
flabel metal2 s 19338 30676 19394 31476 0 FreeSans 224 90 0 0 out[2]
port 28 nsew signal output
flabel metal3 s 28532 25168 29332 25288 0 FreeSans 480 0 0 0 out[30]
port 29 nsew signal output
flabel metal3 s 28532 23808 29332 23928 0 FreeSans 480 0 0 0 out[31]
port 30 nsew signal output
flabel metal3 s 28532 23128 29332 23248 0 FreeSans 480 0 0 0 out[32]
port 31 nsew signal output
flabel metal3 s 28532 22448 29332 22568 0 FreeSans 480 0 0 0 out[33]
port 32 nsew signal output
flabel metal2 s 28354 30676 28410 31476 0 FreeSans 224 90 0 0 out[3]
port 33 nsew signal output
flabel metal2 s 12254 30676 12310 31476 0 FreeSans 224 90 0 0 out[4]
port 34 nsew signal output
flabel metal2 s 18694 30676 18750 31476 0 FreeSans 224 90 0 0 out[5]
port 35 nsew signal output
flabel metal2 s 13542 30676 13598 31476 0 FreeSans 224 90 0 0 out[6]
port 36 nsew signal output
flabel metal2 s 24490 30676 24546 31476 0 FreeSans 224 90 0 0 out[7]
port 37 nsew signal output
flabel metal2 s 20626 30676 20682 31476 0 FreeSans 224 90 0 0 out[8]
port 38 nsew signal output
flabel metal2 s 27710 30676 27766 31476 0 FreeSans 224 90 0 0 out[9]
port 39 nsew signal output
flabel metal2 s 9034 0 9090 800 0 FreeSans 224 90 0 0 prescaler[0]
port 40 nsew signal input
flabel metal3 s 0 23128 800 23248 0 FreeSans 480 0 0 0 prescaler[10]
port 41 nsew signal input
flabel metal3 s 0 22448 800 22568 0 FreeSans 480 0 0 0 prescaler[11]
port 42 nsew signal input
flabel metal3 s 0 23808 800 23928 0 FreeSans 480 0 0 0 prescaler[12]
port 43 nsew signal input
flabel metal3 s 0 21768 800 21888 0 FreeSans 480 0 0 0 prescaler[13]
port 44 nsew signal input
flabel metal2 s 5814 0 5870 800 0 FreeSans 224 90 0 0 prescaler[1]
port 45 nsew signal input
flabel metal3 s 0 11568 800 11688 0 FreeSans 480 0 0 0 prescaler[2]
port 46 nsew signal input
flabel metal3 s 0 13608 800 13728 0 FreeSans 480 0 0 0 prescaler[3]
port 47 nsew signal input
flabel metal3 s 0 14968 800 15088 0 FreeSans 480 0 0 0 prescaler[4]
port 48 nsew signal input
flabel metal3 s 0 17008 800 17128 0 FreeSans 480 0 0 0 prescaler[5]
port 49 nsew signal input
flabel metal3 s 0 19728 800 19848 0 FreeSans 480 0 0 0 prescaler[6]
port 50 nsew signal input
flabel metal3 s 0 21088 800 21208 0 FreeSans 480 0 0 0 prescaler[7]
port 51 nsew signal input
flabel metal3 s 0 20408 800 20528 0 FreeSans 480 0 0 0 prescaler[8]
port 52 nsew signal input
flabel metal3 s 0 19048 800 19168 0 FreeSans 480 0 0 0 prescaler[9]
port 53 nsew signal input
flabel metal3 s 28532 14288 29332 14408 0 FreeSans 480 0 0 0 stop
port 54 nsew signal input
rlabel metal1 14628 28288 14628 28288 0 VGND
rlabel metal1 14628 28832 14628 28832 0 VPWR
rlabel metal1 19205 26962 19205 26962 0 _0000_
rlabel metal2 24058 11084 24058 11084 0 _0001_
rlabel metal1 13202 17850 13202 17850 0 _0002_
rlabel metal1 11914 27064 11914 27064 0 _0003_
rlabel metal1 5704 27438 5704 27438 0 _0004_
rlabel metal1 7866 25262 7866 25262 0 _0005_
rlabel metal1 4048 20910 4048 20910 0 _0006_
rlabel metal1 4600 20026 4600 20026 0 _0007_
rlabel metal1 5244 15470 5244 15470 0 _0008_
rlabel metal2 4922 15776 4922 15776 0 _0009_
rlabel metal1 4600 13906 4600 13906 0 _0010_
rlabel metal2 11638 8704 11638 8704 0 _0011_
rlabel metal1 13570 7344 13570 7344 0 _0012_
rlabel metal2 13846 6766 13846 6766 0 _0013_
rlabel metal2 15318 19686 15318 19686 0 _0014_
rlabel metal1 12650 20400 12650 20400 0 _0015_
rlabel metal1 14444 20910 14444 20910 0 _0016_
rlabel metal1 16698 20468 16698 20468 0 _0017_
rlabel metal1 17894 23528 17894 23528 0 _0018_
rlabel metal1 19090 23120 19090 23120 0 _0019_
rlabel metal1 23598 20774 23598 20774 0 _0020_
rlabel metal1 18584 17510 18584 17510 0 _0021_
rlabel metal1 23690 17612 23690 17612 0 _0022_
rlabel via1 23414 16150 23414 16150 0 _0023_
rlabel metal2 23046 14348 23046 14348 0 _0024_
rlabel metal1 20562 13974 20562 13974 0 _0025_
rlabel metal2 21298 11628 21298 11628 0 _0026_
rlabel metal1 20746 7412 20746 7412 0 _0027_
rlabel metal1 18630 8398 18630 8398 0 _0028_
rlabel metal1 17894 7888 17894 7888 0 _0029_
rlabel metal2 17250 11186 17250 11186 0 _0030_
rlabel metal1 15456 12614 15456 12614 0 _0031_
rlabel metal2 13662 14688 13662 14688 0 _0032_
rlabel metal1 13202 10982 13202 10982 0 _0033_
rlabel via1 12650 9557 12650 9557 0 _0034_
rlabel metal2 13018 6817 13018 6817 0 _0035_
rlabel metal2 16238 7038 16238 7038 0 _0036_
rlabel metal1 24840 10234 24840 10234 0 _0037_
rlabel metal2 23322 7650 23322 7650 0 _0038_
rlabel metal1 22770 26554 22770 26554 0 _0039_
rlabel metal1 22126 26928 22126 26928 0 _0040_
rlabel metal1 26335 24174 26335 24174 0 _0041_
rlabel via1 25798 21862 25798 21862 0 _0042_
rlabel metal2 25622 21658 25622 21658 0 _0043_
rlabel metal1 25635 21658 25635 21658 0 _0044_
rlabel metal1 25024 21386 25024 21386 0 _0045_
rlabel metal2 26174 20910 26174 20910 0 _0046_
rlabel metal1 26128 21658 26128 21658 0 _0047_
rlabel metal2 25806 20876 25806 20876 0 _0048_
rlabel metal1 19596 27438 19596 27438 0 _0049_
rlabel metal2 20470 25568 20470 25568 0 _0050_
rlabel metal1 25208 23834 25208 23834 0 _0051_
rlabel metal2 24242 23290 24242 23290 0 _0052_
rlabel metal1 12972 25874 12972 25874 0 _0053_
rlabel metal1 5566 23188 5566 23188 0 _0054_
rlabel metal2 2530 23902 2530 23902 0 _0055_
rlabel metal1 3450 24140 3450 24140 0 _0056_
rlabel metal2 2530 25806 2530 25806 0 _0057_
rlabel metal1 3634 24208 3634 24208 0 _0058_
rlabel metal2 3634 24548 3634 24548 0 _0059_
rlabel metal1 4508 23290 4508 23290 0 _0060_
rlabel metal1 4554 24106 4554 24106 0 _0061_
rlabel metal2 5198 24378 5198 24378 0 _0062_
rlabel metal1 4002 26996 4002 26996 0 _0063_
rlabel metal1 2622 26928 2622 26928 0 _0064_
rlabel metal1 3680 26350 3680 26350 0 _0065_
rlabel metal1 3542 26894 3542 26894 0 _0066_
rlabel metal1 3956 26554 3956 26554 0 _0067_
rlabel metal1 4876 24174 4876 24174 0 _0068_
rlabel metal1 5244 23154 5244 23154 0 _0069_
rlabel metal2 5658 22814 5658 22814 0 _0070_
rlabel metal1 6026 23086 6026 23086 0 _0071_
rlabel metal1 4738 26894 4738 26894 0 _0072_
rlabel metal2 5428 26894 5428 26894 0 _0073_
rlabel metal2 6118 27438 6118 27438 0 _0074_
rlabel metal2 5566 27132 5566 27132 0 _0075_
rlabel metal1 5152 26554 5152 26554 0 _0076_
rlabel metal1 5553 27098 5553 27098 0 _0077_
rlabel metal1 5566 26826 5566 26826 0 _0078_
rlabel metal1 5658 26384 5658 26384 0 _0079_
rlabel metal2 6302 24684 6302 24684 0 _0080_
rlabel metal1 7176 22678 7176 22678 0 _0081_
rlabel metal2 7314 21726 7314 21726 0 _0082_
rlabel metal1 7682 22406 7682 22406 0 _0083_
rlabel metal1 6118 25262 6118 25262 0 _0084_
rlabel metal1 6532 26418 6532 26418 0 _0085_
rlabel metal2 6578 25772 6578 25772 0 _0086_
rlabel metal1 7682 24786 7682 24786 0 _0087_
rlabel metal1 7360 24174 7360 24174 0 _0088_
rlabel metal2 8142 24582 8142 24582 0 _0089_
rlabel metal1 8050 23018 8050 23018 0 _0090_
rlabel metal2 8878 22950 8878 22950 0 _0091_
rlabel metal1 10626 23120 10626 23120 0 _0092_
rlabel metal1 8694 22712 8694 22712 0 _0093_
rlabel metal1 9614 22984 9614 22984 0 _0094_
rlabel metal1 5014 11186 5014 11186 0 _0095_
rlabel metal2 2714 10302 2714 10302 0 _0096_
rlabel metal1 2714 10676 2714 10676 0 _0097_
rlabel metal1 9568 11118 9568 11118 0 _0098_
rlabel metal2 4646 13498 4646 13498 0 _0099_
rlabel metal2 2438 12546 2438 12546 0 _0100_
rlabel metal1 2254 13838 2254 13838 0 _0101_
rlabel metal1 2944 11118 2944 11118 0 _0102_
rlabel metal1 3496 11186 3496 11186 0 _0103_
rlabel metal1 4002 9996 4002 9996 0 _0104_
rlabel metal2 4094 10268 4094 10268 0 _0105_
rlabel metal2 4554 11798 4554 11798 0 _0106_
rlabel metal1 2898 13260 2898 13260 0 _0107_
rlabel metal1 4462 15436 4462 15436 0 _0108_
rlabel metal1 2208 16626 2208 16626 0 _0109_
rlabel metal1 2254 17068 2254 17068 0 _0110_
rlabel metal2 2346 14858 2346 14858 0 _0111_
rlabel metal1 3542 13838 3542 13838 0 _0112_
rlabel metal2 2990 13600 2990 13600 0 _0113_
rlabel metal1 3542 13158 3542 13158 0 _0114_
rlabel metal1 4646 11696 4646 11696 0 _0115_
rlabel metal1 4830 11730 4830 11730 0 _0116_
rlabel metal1 4968 12818 4968 12818 0 _0117_
rlabel metal2 2806 14212 2806 14212 0 _0118_
rlabel metal1 2852 15130 2852 15130 0 _0119_
rlabel metal1 5014 18292 5014 18292 0 _0120_
rlabel metal1 2024 19822 2024 19822 0 _0121_
rlabel metal1 2438 19856 2438 19856 0 _0122_
rlabel metal1 2622 17245 2622 17245 0 _0123_
rlabel metal2 2990 16762 2990 16762 0 _0124_
rlabel metal2 3266 16932 3266 16932 0 _0125_
rlabel metal2 3266 14858 3266 14858 0 _0126_
rlabel metal2 3634 14212 3634 14212 0 _0127_
rlabel metal1 4370 14518 4370 14518 0 _0128_
rlabel metal1 5382 12893 5382 12893 0 _0129_
rlabel metal1 7360 13226 7360 13226 0 _0130_
rlabel metal1 6167 12206 6167 12206 0 _0131_
rlabel metal1 7130 13294 7130 13294 0 _0132_
rlabel metal2 5474 14654 5474 14654 0 _0133_
rlabel metal2 3542 18428 3542 18428 0 _0134_
rlabel metal1 5520 20366 5520 20366 0 _0135_
rlabel metal1 1978 21624 1978 21624 0 _0136_
rlabel metal1 2944 22542 2944 22542 0 _0137_
rlabel metal2 2898 20842 2898 20842 0 _0138_
rlabel metal1 3220 19278 3220 19278 0 _0139_
rlabel metal2 3726 18768 3726 18768 0 _0140_
rlabel metal2 4002 17680 4002 17680 0 _0141_
rlabel metal1 3772 16626 3772 16626 0 _0142_
rlabel metal2 3910 16524 3910 16524 0 _0143_
rlabel metal2 4646 16252 4646 16252 0 _0144_
rlabel metal1 4968 14382 4968 14382 0 _0145_
rlabel metal2 6210 14586 6210 14586 0 _0146_
rlabel metal1 6578 14450 6578 14450 0 _0147_
rlabel metal1 6946 13838 6946 13838 0 _0148_
rlabel metal1 8326 13328 8326 13328 0 _0149_
rlabel metal1 6578 8500 6578 8500 0 _0150_
rlabel metal1 5244 7174 5244 7174 0 _0151_
rlabel metal2 4830 7684 4830 7684 0 _0152_
rlabel metal1 4370 7888 4370 7888 0 _0153_
rlabel metal1 5750 7820 5750 7820 0 _0154_
rlabel metal1 5750 7344 5750 7344 0 _0155_
rlabel metal2 5474 7582 5474 7582 0 _0156_
rlabel metal2 5382 8704 5382 8704 0 _0157_
rlabel metal1 4922 9010 4922 9010 0 _0158_
rlabel metal1 5612 8602 5612 8602 0 _0159_
rlabel metal2 5934 8670 5934 8670 0 _0160_
rlabel metal1 6486 10642 6486 10642 0 _0161_
rlabel metal2 6486 10778 6486 10778 0 _0162_
rlabel metal2 5842 10914 5842 10914 0 _0163_
rlabel metal1 7544 10574 7544 10574 0 _0164_
rlabel metal1 7498 12750 7498 12750 0 _0165_
rlabel metal1 7537 12818 7537 12818 0 _0166_
rlabel metal2 8280 13294 8280 13294 0 _0167_
rlabel metal1 9522 12818 9522 12818 0 _0168_
rlabel metal1 8924 10098 8924 10098 0 _0169_
rlabel metal2 7590 7004 7590 7004 0 _0170_
rlabel metal1 7038 6290 7038 6290 0 _0171_
rlabel metal2 8694 10880 8694 10880 0 _0172_
rlabel metal1 8602 7514 8602 7514 0 _0173_
rlabel metal2 8786 6460 8786 6460 0 _0174_
rlabel metal2 8694 6154 8694 6154 0 _0175_
rlabel metal1 9614 6290 9614 6290 0 _0176_
rlabel metal1 8648 6222 8648 6222 0 _0177_
rlabel metal2 8510 6290 8510 6290 0 _0178_
rlabel metal2 8050 7174 8050 7174 0 _0179_
rlabel metal2 8418 7106 8418 7106 0 _0180_
rlabel metal2 8050 7990 8050 7990 0 _0181_
rlabel metal1 7958 8364 7958 8364 0 _0182_
rlabel metal2 8970 9248 8970 9248 0 _0183_
rlabel metal1 8970 8534 8970 8534 0 _0184_
rlabel metal2 9154 7174 9154 7174 0 _0185_
rlabel metal1 9660 6766 9660 6766 0 _0186_
rlabel metal1 7682 9996 7682 9996 0 _0187_
rlabel metal1 8740 10574 8740 10574 0 _0188_
rlabel metal1 9614 11696 9614 11696 0 _0189_
rlabel metal1 9890 10710 9890 10710 0 _0190_
rlabel metal1 9246 7344 9246 7344 0 _0191_
rlabel metal1 10074 7718 10074 7718 0 _0192_
rlabel metal1 9798 8908 9798 8908 0 _0193_
rlabel metal1 9614 12750 9614 12750 0 _0194_
rlabel metal2 9246 13498 9246 13498 0 _0195_
rlabel metal1 8234 13770 8234 13770 0 _0196_
rlabel metal2 8786 14484 8786 14484 0 _0197_
rlabel metal1 8786 15606 8786 15606 0 _0198_
rlabel metal2 8418 14756 8418 14756 0 _0199_
rlabel metal1 5106 16592 5106 16592 0 _0200_
rlabel metal1 4462 19380 4462 19380 0 _0201_
rlabel metal2 3818 21318 3818 21318 0 _0202_
rlabel metal2 3082 23120 3082 23120 0 _0203_
rlabel metal2 3910 22236 3910 22236 0 _0204_
rlabel metal1 4186 21964 4186 21964 0 _0205_
rlabel metal2 4738 20502 4738 20502 0 _0206_
rlabel metal2 5566 19108 5566 19108 0 _0207_
rlabel metal2 5290 18496 5290 18496 0 _0208_
rlabel metal1 5934 16558 5934 16558 0 _0209_
rlabel metal1 5428 16422 5428 16422 0 _0210_
rlabel metal2 6946 16354 6946 16354 0 _0211_
rlabel metal1 8188 15538 8188 15538 0 _0212_
rlabel metal1 8740 16150 8740 16150 0 _0213_
rlabel metal2 9890 15266 9890 15266 0 _0214_
rlabel metal1 5750 18768 5750 18768 0 _0215_
rlabel metal2 4646 21692 4646 21692 0 _0216_
rlabel metal2 5014 21216 5014 21216 0 _0217_
rlabel metal1 5106 20774 5106 20774 0 _0218_
rlabel metal2 5750 20672 5750 20672 0 _0219_
rlabel metal2 6486 19550 6486 19550 0 _0220_
rlabel metal1 6670 18190 6670 18190 0 _0221_
rlabel metal1 7636 18190 7636 18190 0 _0222_
rlabel metal2 8602 17374 8602 17374 0 _0223_
rlabel metal2 8050 16864 8050 16864 0 _0224_
rlabel metal1 9338 16592 9338 16592 0 _0225_
rlabel metal2 9430 17476 9430 17476 0 _0226_
rlabel metal1 6210 20910 6210 20910 0 _0227_
rlabel metal1 6808 20910 6808 20910 0 _0228_
rlabel metal2 7130 20638 7130 20638 0 _0229_
rlabel metal2 7774 20672 7774 20672 0 _0230_
rlabel metal2 7866 19516 7866 19516 0 _0231_
rlabel metal2 7958 18768 7958 18768 0 _0232_
rlabel metal2 10994 18258 10994 18258 0 _0233_
rlabel metal2 9706 18938 9706 18938 0 _0234_
rlabel metal1 10028 17170 10028 17170 0 _0235_
rlabel metal1 8326 19346 8326 19346 0 _0236_
rlabel metal2 8142 20400 8142 20400 0 _0237_
rlabel metal1 10120 18734 10120 18734 0 _0238_
rlabel metal1 10212 18598 10212 18598 0 _0239_
rlabel metal2 7590 16082 7590 16082 0 _0240_
rlabel metal1 8510 18190 8510 18190 0 _0241_
rlabel metal2 9430 20468 9430 20468 0 _0242_
rlabel metal2 8234 18938 8234 18938 0 _0243_
rlabel via1 8329 18598 8329 18598 0 _0244_
rlabel metal2 9246 19856 9246 19856 0 _0245_
rlabel metal1 9522 22066 9522 22066 0 _0246_
rlabel metal1 9982 24174 9982 24174 0 _0247_
rlabel metal1 6854 27506 6854 27506 0 _0248_
rlabel metal1 6992 26962 6992 26962 0 _0249_
rlabel metal2 7682 26554 7682 26554 0 _0250_
rlabel metal1 7498 26384 7498 26384 0 _0251_
rlabel metal1 7728 25942 7728 25942 0 _0252_
rlabel metal1 8602 26384 8602 26384 0 _0253_
rlabel metal1 8050 25296 8050 25296 0 _0254_
rlabel metal2 8418 24956 8418 24956 0 _0255_
rlabel metal1 8878 24174 8878 24174 0 _0256_
rlabel via1 9425 24174 9425 24174 0 _0257_
rlabel metal1 9384 23086 9384 23086 0 _0258_
rlabel metal1 11224 27438 11224 27438 0 _0259_
rlabel metal1 10810 27404 10810 27404 0 _0260_
rlabel metal2 12006 27166 12006 27166 0 _0261_
rlabel metal2 10534 26962 10534 26962 0 _0262_
rlabel metal1 10626 26418 10626 26418 0 _0263_
rlabel metal1 10258 26860 10258 26860 0 _0264_
rlabel metal1 12282 24820 12282 24820 0 _0265_
rlabel metal1 11132 26554 11132 26554 0 _0266_
rlabel metal1 9798 26860 9798 26860 0 _0267_
rlabel metal2 9798 26554 9798 26554 0 _0268_
rlabel metal1 10626 25908 10626 25908 0 _0269_
rlabel metal2 10442 26044 10442 26044 0 _0270_
rlabel metal1 15134 25364 15134 25364 0 _0271_
rlabel metal2 8786 26554 8786 26554 0 _0272_
rlabel metal1 15502 25228 15502 25228 0 _0273_
rlabel metal1 9016 25262 9016 25262 0 _0274_
rlabel metal1 9706 24786 9706 24786 0 _0275_
rlabel metal1 10120 24582 10120 24582 0 _0276_
rlabel metal1 9844 23086 9844 23086 0 _0277_
rlabel metal2 11822 23698 11822 23698 0 _0278_
rlabel metal1 9660 23766 9660 23766 0 _0279_
rlabel metal2 10442 24004 10442 24004 0 _0280_
rlabel metal2 10534 24956 10534 24956 0 _0281_
rlabel metal1 11316 24718 11316 24718 0 _0282_
rlabel metal2 12558 26044 12558 26044 0 _0283_
rlabel metal1 12650 26350 12650 26350 0 _0284_
rlabel metal1 12420 26962 12420 26962 0 _0285_
rlabel metal2 12558 26656 12558 26656 0 _0286_
rlabel metal1 12144 24786 12144 24786 0 _0287_
rlabel metal1 12190 25262 12190 25262 0 _0288_
rlabel metal1 12926 23494 12926 23494 0 _0289_
rlabel metal1 12098 23766 12098 23766 0 _0290_
rlabel metal2 14582 20128 14582 20128 0 _0291_
rlabel metal1 14858 18292 14858 18292 0 _0292_
rlabel metal1 14858 18054 14858 18054 0 _0293_
rlabel metal1 15502 20910 15502 20910 0 _0294_
rlabel metal1 14766 20026 14766 20026 0 _0295_
rlabel metal2 16238 21216 16238 21216 0 _0296_
rlabel metal1 16330 21964 16330 21964 0 _0297_
rlabel metal2 12926 24106 12926 24106 0 _0298_
rlabel metal1 12144 16558 12144 16558 0 _0299_
rlabel metal1 14030 21522 14030 21522 0 _0300_
rlabel metal1 14628 22066 14628 22066 0 _0301_
rlabel metal2 13202 24582 13202 24582 0 _0302_
rlabel metal1 16284 14926 16284 14926 0 _0303_
rlabel metal1 13992 22746 13992 22746 0 _0304_
rlabel metal1 16468 21862 16468 21862 0 _0305_
rlabel metal1 17618 21488 17618 21488 0 _0306_
rlabel metal1 18308 16014 18308 16014 0 _0307_
rlabel metal1 14122 24140 14122 24140 0 _0308_
rlabel metal2 15962 24140 15962 24140 0 _0309_
rlabel metal2 15778 24140 15778 24140 0 _0310_
rlabel metal2 16790 24956 16790 24956 0 _0311_
rlabel metal2 16698 24990 16698 24990 0 _0312_
rlabel metal1 15916 23494 15916 23494 0 _0313_
rlabel metal1 17434 23698 17434 23698 0 _0314_
rlabel metal2 17802 24378 17802 24378 0 _0315_
rlabel metal1 17434 23834 17434 23834 0 _0316_
rlabel metal1 14306 24242 14306 24242 0 _0317_
rlabel metal1 19044 19890 19044 19890 0 _0318_
rlabel metal1 17948 23834 17948 23834 0 _0319_
rlabel metal2 18078 21148 18078 21148 0 _0320_
rlabel metal1 18722 23154 18722 23154 0 _0321_
rlabel metal1 16054 23086 16054 23086 0 _0322_
rlabel metal1 19504 19346 19504 19346 0 _0323_
rlabel metal1 19734 23222 19734 23222 0 _0324_
rlabel metal1 19366 23290 19366 23290 0 _0325_
rlabel metal2 21574 20400 21574 20400 0 _0326_
rlabel metal2 20470 22882 20470 22882 0 _0327_
rlabel metal1 18262 23630 18262 23630 0 _0328_
rlabel metal1 17434 23562 17434 23562 0 _0329_
rlabel metal1 16974 22066 16974 22066 0 _0330_
rlabel metal2 17158 21692 17158 21692 0 _0331_
rlabel metal2 14490 21828 14490 21828 0 _0332_
rlabel metal2 15226 21420 15226 21420 0 _0333_
rlabel metal2 15134 20366 15134 20366 0 _0334_
rlabel via2 22494 19363 22494 19363 0 _0335_
rlabel metal2 15502 20434 15502 20434 0 _0336_
rlabel metal2 20838 22916 20838 22916 0 _0337_
rlabel metal1 19964 23018 19964 23018 0 _0338_
rlabel metal1 17710 21012 17710 21012 0 _0339_
rlabel metal1 17940 15946 17940 15946 0 _0340_
rlabel metal2 9890 17612 9890 17612 0 _0341_
rlabel metal1 11040 17850 11040 17850 0 _0342_
rlabel metal1 18860 17646 18860 17646 0 _0343_
rlabel metal1 17664 16558 17664 16558 0 _0344_
rlabel metal1 15916 17170 15916 17170 0 _0345_
rlabel metal2 20746 17068 20746 17068 0 _0346_
rlabel metal1 21022 16524 21022 16524 0 _0347_
rlabel metal1 21068 16014 21068 16014 0 _0348_
rlabel metal1 9200 15946 9200 15946 0 _0349_
rlabel metal2 22126 13022 22126 13022 0 _0350_
rlabel metal1 17066 17306 17066 17306 0 _0351_
rlabel metal2 21390 15742 21390 15742 0 _0352_
rlabel metal1 21574 15436 21574 15436 0 _0353_
rlabel via1 21482 14926 21482 14926 0 _0354_
rlabel metal1 20792 15130 20792 15130 0 _0355_
rlabel metal1 19642 15572 19642 15572 0 _0356_
rlabel metal2 9154 13532 9154 13532 0 _0357_
rlabel metal2 19826 13396 19826 13396 0 _0358_
rlabel metal1 18630 13872 18630 13872 0 _0359_
rlabel metal1 20286 11594 20286 11594 0 _0360_
rlabel metal1 20838 11730 20838 11730 0 _0361_
rlabel metal2 19642 12240 19642 12240 0 _0362_
rlabel metal1 18262 12954 18262 12954 0 _0363_
rlabel metal1 20056 11594 20056 11594 0 _0364_
rlabel metal1 19412 14790 19412 14790 0 _0365_
rlabel metal1 9936 7446 9936 7446 0 _0366_
rlabel via1 15985 7854 15985 7854 0 _0367_
rlabel metal1 16836 10234 16836 10234 0 _0368_
rlabel metal1 9936 7378 9936 7378 0 _0369_
rlabel metal1 16192 10030 16192 10030 0 _0370_
rlabel metal1 17066 10506 17066 10506 0 _0371_
rlabel metal1 9476 10642 9476 10642 0 _0372_
rlabel metal1 14168 11730 14168 11730 0 _0373_
rlabel metal1 15548 14382 15548 14382 0 _0374_
rlabel metal1 16192 10982 16192 10982 0 _0375_
rlabel metal1 9292 11730 9292 11730 0 _0376_
rlabel metal2 12558 13209 12558 13209 0 _0377_
rlabel metal2 14490 11084 14490 11084 0 _0378_
rlabel metal1 13708 8942 13708 8942 0 _0379_
rlabel metal1 13708 8534 13708 8534 0 _0380_
rlabel metal1 12972 9146 12972 9146 0 _0381_
rlabel metal2 14030 10846 14030 10846 0 _0382_
rlabel metal1 12052 10234 12052 10234 0 _0383_
rlabel metal2 11822 10914 11822 10914 0 _0384_
rlabel metal1 13110 10574 13110 10574 0 _0385_
rlabel metal2 12650 10812 12650 10812 0 _0386_
rlabel metal1 14214 10608 14214 10608 0 _0387_
rlabel viali 16971 10574 16971 10574 0 _0388_
rlabel metal1 17986 10710 17986 10710 0 _0389_
rlabel metal1 9384 9690 9384 9690 0 _0390_
rlabel metal2 19642 9656 19642 9656 0 _0391_
rlabel metal2 20654 8058 20654 8058 0 _0392_
rlabel metal1 19228 10098 19228 10098 0 _0393_
rlabel metal1 18998 9962 18998 9962 0 _0394_
rlabel metal2 9706 8772 9706 8772 0 _0395_
rlabel metal1 18170 13974 18170 13974 0 _0396_
rlabel metal1 18676 9690 18676 9690 0 _0397_
rlabel metal1 18446 14926 18446 14926 0 _0398_
rlabel metal1 19136 11186 19136 11186 0 _0399_
rlabel metal2 18998 10234 18998 10234 0 _0400_
rlabel metal2 19826 11764 19826 11764 0 _0401_
rlabel metal1 19366 12410 19366 12410 0 _0402_
rlabel metal1 21298 17068 21298 17068 0 _0403_
rlabel metal2 20838 16524 20838 16524 0 _0404_
rlabel metal2 21114 15776 21114 15776 0 _0405_
rlabel metal2 19826 15674 19826 15674 0 _0406_
rlabel metal1 18998 21488 18998 21488 0 _0407_
rlabel metal2 22586 14994 22586 14994 0 _0408_
rlabel metal1 18124 21114 18124 21114 0 _0409_
rlabel metal1 23322 19142 23322 19142 0 _0410_
rlabel metal1 23966 10506 23966 10506 0 _0411_
rlabel metal1 14766 8534 14766 8534 0 _0412_
rlabel metal1 14306 8602 14306 8602 0 _0413_
rlabel metal2 14766 10438 14766 10438 0 _0414_
rlabel via2 17526 10659 17526 10659 0 _0415_
rlabel metal1 18308 14994 18308 14994 0 _0416_
rlabel metal1 18722 15130 18722 15130 0 _0417_
rlabel metal1 22954 15402 22954 15402 0 _0418_
rlabel metal1 23782 17102 23782 17102 0 _0419_
rlabel metal1 10212 11050 10212 11050 0 _0420_
rlabel metal1 10718 11322 10718 11322 0 _0421_
rlabel metal2 20102 12257 20102 12257 0 _0422_
rlabel metal1 22494 12750 22494 12750 0 _0423_
rlabel metal1 23690 12716 23690 12716 0 _0424_
rlabel metal1 24104 12886 24104 12886 0 _0425_
rlabel metal1 22862 13498 22862 13498 0 _0426_
rlabel metal1 23782 11220 23782 11220 0 _0427_
rlabel metal1 24472 10438 24472 10438 0 _0428_
rlabel metal1 24204 10778 24204 10778 0 _0429_
rlabel metal2 23690 9146 23690 9146 0 _0430_
rlabel metal2 23414 8772 23414 8772 0 _0431_
rlabel metal1 23598 8364 23598 8364 0 _0432_
rlabel metal1 23598 8976 23598 8976 0 _0433_
rlabel metal2 23782 8466 23782 8466 0 _0434_
rlabel metal2 14214 7259 14214 7259 0 _0435_
rlabel metal2 22034 24514 22034 24514 0 _0436_
rlabel metal1 21850 24786 21850 24786 0 _0437_
rlabel metal1 23552 23698 23552 23698 0 _0438_
rlabel metal2 21574 24004 21574 24004 0 _0439_
rlabel metal1 22724 23086 22724 23086 0 _0440_
rlabel metal2 15226 7582 15226 7582 0 _0441_
rlabel metal1 14766 6766 14766 6766 0 _0442_
rlabel metal2 15134 7174 15134 7174 0 _0443_
rlabel metal1 15456 7378 15456 7378 0 _0444_
rlabel metal1 12696 6970 12696 6970 0 _0445_
rlabel metal2 13386 7548 13386 7548 0 _0446_
rlabel metal2 13110 7072 13110 7072 0 _0447_
rlabel metal1 12880 7514 12880 7514 0 _0448_
rlabel metal1 12926 6630 12926 6630 0 _0449_
rlabel metal2 12282 9146 12282 9146 0 _0450_
rlabel metal1 13064 9554 13064 9554 0 _0451_
rlabel metal1 13248 9418 13248 9418 0 _0452_
rlabel metal2 12374 9146 12374 9146 0 _0453_
rlabel metal2 12098 9486 12098 9486 0 _0454_
rlabel metal1 12466 8976 12466 8976 0 _0455_
rlabel metal1 12604 11866 12604 11866 0 _0456_
rlabel metal1 13156 10234 13156 10234 0 _0457_
rlabel metal1 12558 11050 12558 11050 0 _0458_
rlabel metal1 12650 11322 12650 11322 0 _0459_
rlabel metal2 13202 12036 13202 12036 0 _0460_
rlabel metal1 12466 16490 12466 16490 0 _0461_
rlabel metal1 12880 14586 12880 14586 0 _0462_
rlabel metal1 14904 13294 14904 13294 0 _0463_
rlabel metal2 13846 13600 13846 13600 0 _0464_
rlabel metal2 13478 14416 13478 14416 0 _0465_
rlabel metal1 16100 12954 16100 12954 0 _0466_
rlabel metal1 15916 13226 15916 13226 0 _0467_
rlabel metal1 16054 13328 16054 13328 0 _0468_
rlabel metal1 15226 14382 15226 14382 0 _0469_
rlabel metal2 14858 13940 14858 13940 0 _0470_
rlabel metal1 17342 11798 17342 11798 0 _0471_
rlabel metal1 16054 12308 16054 12308 0 _0472_
rlabel metal1 15732 11322 15732 11322 0 _0473_
rlabel metal2 15962 11900 15962 11900 0 _0474_
rlabel metal2 16330 11407 16330 11407 0 _0475_
rlabel metal1 16974 7378 16974 7378 0 _0476_
rlabel metal2 17158 8636 17158 8636 0 _0477_
rlabel metal2 17342 8806 17342 8806 0 _0478_
rlabel metal2 16790 7820 16790 7820 0 _0479_
rlabel metal1 17296 7378 17296 7378 0 _0480_
rlabel metal2 19090 7548 19090 7548 0 _0481_
rlabel metal2 20194 9792 20194 9792 0 _0482_
rlabel metal1 19780 8058 19780 8058 0 _0483_
rlabel metal2 19274 7514 19274 7514 0 _0484_
rlabel metal1 20884 7242 20884 7242 0 _0485_
rlabel metal1 22218 7412 22218 7412 0 _0486_
rlabel metal2 21666 7582 21666 7582 0 _0487_
rlabel metal1 20608 7514 20608 7514 0 _0488_
rlabel metal1 20930 10710 20930 10710 0 _0489_
rlabel metal1 21574 13260 21574 13260 0 _0490_
rlabel metal2 22218 9894 22218 9894 0 _0491_
rlabel metal2 21850 10132 21850 10132 0 _0492_
rlabel metal1 20700 10642 20700 10642 0 _0493_
rlabel metal2 19550 13158 19550 13158 0 _0494_
rlabel metal1 21942 13974 21942 13974 0 _0495_
rlabel metal1 21620 13498 21620 13498 0 _0496_
rlabel metal1 20746 13872 20746 13872 0 _0497_
rlabel metal1 19458 13328 19458 13328 0 _0498_
rlabel via1 19642 13498 19642 13498 0 _0499_
rlabel metal1 23414 13940 23414 13940 0 _0500_
rlabel metal1 24886 13430 24886 13430 0 _0501_
rlabel metal1 24012 13498 24012 13498 0 _0502_
rlabel metal1 23000 16218 23000 16218 0 _0503_
rlabel metal1 24610 17170 24610 17170 0 _0504_
rlabel metal1 24380 15606 24380 15606 0 _0505_
rlabel metal1 23552 15674 23552 15674 0 _0506_
rlabel metal1 23322 15980 23322 15980 0 _0507_
rlabel metal2 22126 16286 22126 16286 0 _0508_
rlabel metal1 24242 17136 24242 17136 0 _0509_
rlabel metal2 24426 17374 24426 17374 0 _0510_
rlabel metal1 23414 17204 23414 17204 0 _0511_
rlabel metal1 24104 17306 24104 17306 0 _0512_
rlabel metal1 22448 17782 22448 17782 0 _0513_
rlabel metal1 18032 16762 18032 16762 0 _0514_
rlabel metal1 17894 17680 17894 17680 0 _0515_
rlabel metal1 21988 20230 21988 20230 0 _0516_
rlabel metal2 23414 20468 23414 20468 0 _0517_
rlabel metal1 23548 19482 23548 19482 0 _0518_
rlabel via1 22042 20570 22042 20570 0 _0519_
rlabel metal2 22218 20672 22218 20672 0 _0520_
rlabel metal2 22494 20400 22494 20400 0 _0521_
rlabel metal1 20700 20910 20700 20910 0 _0522_
rlabel metal1 21068 20842 21068 20842 0 _0523_
rlabel metal2 20378 20332 20378 20332 0 _0524_
rlabel metal2 20194 20434 20194 20434 0 _0525_
rlabel metal2 20102 20570 20102 20570 0 _0526_
rlabel metal2 18538 19856 18538 19856 0 _0527_
rlabel metal2 19642 21726 19642 21726 0 _0528_
rlabel metal1 18446 19380 18446 19380 0 _0529_
rlabel metal2 18722 20060 18722 20060 0 _0530_
rlabel metal2 18906 16558 18906 16558 0 _0531_
rlabel metal2 17342 22372 17342 22372 0 _0532_
rlabel metal1 17204 21998 17204 21998 0 _0533_
rlabel metal1 17618 21862 17618 21862 0 _0534_
rlabel metal1 16744 20366 16744 20366 0 _0535_
rlabel metal1 16422 20026 16422 20026 0 _0536_
rlabel metal1 13064 20570 13064 20570 0 _0537_
rlabel via1 13386 19227 13386 19227 0 _0538_
rlabel metal1 13064 21590 13064 21590 0 _0539_
rlabel metal2 13018 21148 13018 21148 0 _0540_
rlabel metal1 13708 20910 13708 20910 0 _0541_
rlabel metal1 15778 14790 15778 14790 0 _0542_
rlabel metal1 12420 20434 12420 20434 0 _0543_
rlabel metal1 12834 19720 12834 19720 0 _0544_
rlabel metal1 13064 19822 13064 19822 0 _0545_
rlabel metal2 12374 20196 12374 20196 0 _0546_
rlabel metal1 15548 18258 15548 18258 0 _0547_
rlabel metal1 15686 18054 15686 18054 0 _0548_
rlabel metal1 16100 18122 16100 18122 0 _0549_
rlabel metal2 12926 16762 12926 16762 0 _0550_
rlabel metal2 13202 18768 13202 18768 0 _0551_
rlabel metal2 13294 18428 13294 18428 0 _0552_
rlabel metal1 12834 16626 12834 16626 0 _0553_
rlabel metal2 23414 10982 23414 10982 0 _0554_
rlabel metal1 22908 12886 22908 12886 0 _0555_
rlabel metal2 23230 12988 23230 12988 0 _0556_
rlabel metal1 23460 12750 23460 12750 0 _0557_
rlabel metal1 23460 12614 23460 12614 0 _0558_
rlabel metal1 17296 14042 17296 14042 0 _0559_
rlabel metal1 16376 8058 16376 8058 0 _0560_
rlabel metal1 17802 7514 17802 7514 0 _0561_
rlabel metal2 16606 7667 16606 7667 0 _0562_
rlabel metal2 19826 12716 19826 12716 0 _0563_
rlabel metal1 20746 17714 20746 17714 0 _0564_
rlabel metal2 21390 17000 21390 17000 0 _0565_
rlabel metal1 20056 17714 20056 17714 0 _0566_
rlabel metal2 20286 17340 20286 17340 0 _0567_
rlabel metal1 16192 16966 16192 16966 0 _0568_
rlabel metal1 15318 17170 15318 17170 0 _0569_
rlabel metal1 15640 14586 15640 14586 0 _0570_
rlabel metal1 19688 17238 19688 17238 0 _0571_
rlabel metal2 21850 17255 21850 17255 0 _0572_
rlabel metal1 18630 13396 18630 13396 0 _0573_
rlabel metal1 15134 13430 15134 13430 0 _0574_
rlabel metal1 17204 14450 17204 14450 0 _0575_
rlabel metal1 17204 17170 17204 17170 0 _0576_
rlabel metal2 15410 14484 15410 14484 0 _0577_
rlabel metal2 22264 19686 22264 19686 0 _0578_
rlabel metal2 15226 13673 15226 13673 0 _0579_
rlabel metal2 14858 16048 14858 16048 0 _0580_
rlabel metal1 15594 17034 15594 17034 0 _0581_
rlabel metal1 13202 13294 13202 13294 0 _0582_
rlabel metal1 16790 16966 16790 16966 0 _0583_
rlabel metal1 13064 16082 13064 16082 0 _0584_
rlabel metal2 12834 15504 12834 15504 0 _0585_
rlabel metal1 14950 16014 14950 16014 0 _0586_
rlabel metal2 12834 16286 12834 16286 0 _0587_
rlabel metal1 15180 15946 15180 15946 0 _0588_
rlabel metal3 18653 16524 18653 16524 0 _0589_
rlabel metal1 17986 16082 17986 16082 0 _0590_
rlabel metal2 18170 17782 18170 17782 0 _0591_
rlabel metal2 17986 14926 17986 14926 0 _0592_
rlabel metal1 14996 7514 14996 7514 0 _0593_
rlabel metal1 15456 14314 15456 14314 0 _0594_
rlabel metal1 17342 16218 17342 16218 0 _0595_
rlabel metal1 22034 17136 22034 17136 0 _0596_
rlabel metal1 27094 25194 27094 25194 0 _0597_
rlabel metal2 25622 24344 25622 24344 0 _0598_
rlabel metal1 26772 25194 26772 25194 0 _0599_
rlabel metal1 26726 25942 26726 25942 0 _0600_
rlabel metal1 27186 24718 27186 24718 0 _0601_
rlabel metal1 18630 26928 18630 26928 0 _0602_
rlabel metal2 26358 25330 26358 25330 0 _0603_
rlabel metal2 26450 25432 26450 25432 0 _0604_
rlabel metal2 18722 28220 18722 28220 0 _0605_
rlabel metal1 19366 27438 19366 27438 0 _0606_
rlabel metal1 27002 27404 27002 27404 0 _0607_
rlabel metal2 18354 26656 18354 26656 0 _0608_
rlabel metal1 17250 27472 17250 27472 0 _0609_
rlabel metal1 20378 26996 20378 26996 0 _0610_
rlabel metal2 21114 27778 21114 27778 0 _0611_
rlabel metal2 22126 27676 22126 27676 0 _0612_
rlabel metal1 24518 27098 24518 27098 0 _0613_
rlabel metal1 20010 27098 20010 27098 0 _0614_
rlabel metal1 26036 26962 26036 26962 0 _0615_
rlabel metal2 21022 27506 21022 27506 0 _0616_
rlabel metal1 25116 27642 25116 27642 0 _0617_
rlabel metal1 17940 26962 17940 26962 0 _0618_
rlabel metal1 19182 27982 19182 27982 0 _0619_
rlabel metal1 26136 26010 26136 26010 0 _0620_
rlabel via3 20539 15300 20539 15300 0 clk
rlabel metal1 24748 11730 24748 11730 0 clk_divider.count_out\[0\]
rlabel metal2 15410 11628 15410 11628 0 clk_divider.count_out\[10\]
rlabel metal1 18170 7344 18170 7344 0 clk_divider.count_out\[11\]
rlabel metal2 18998 7650 18998 7650 0 clk_divider.count_out\[12\]
rlabel metal1 21252 7854 21252 7854 0 clk_divider.count_out\[13\]
rlabel metal1 20654 9962 20654 9962 0 clk_divider.count_out\[14\]
rlabel metal1 21436 13498 21436 13498 0 clk_divider.count_out\[15\]
rlabel metal2 24610 14212 24610 14212 0 clk_divider.count_out\[16\]
rlabel metal1 21712 15470 21712 15470 0 clk_divider.count_out\[17\]
rlabel metal1 22586 17680 22586 17680 0 clk_divider.count_out\[18\]
rlabel metal2 23414 19635 23414 19635 0 clk_divider.count_out\[19\]
rlabel metal1 24978 9962 24978 9962 0 clk_divider.count_out\[1\]
rlabel metal2 24058 19550 24058 19550 0 clk_divider.count_out\[20\]
rlabel metal2 21114 21216 21114 21216 0 clk_divider.count_out\[21\]
rlabel metal2 18630 24038 18630 24038 0 clk_divider.count_out\[22\]
rlabel metal1 16790 22644 16790 22644 0 clk_divider.count_out\[23\]
rlabel metal1 12512 21522 12512 21522 0 clk_divider.count_out\[24\]
rlabel metal1 13340 19822 13340 19822 0 clk_divider.count_out\[25\]
rlabel metal2 15778 18292 15778 18292 0 clk_divider.count_out\[26\]
rlabel metal1 13662 16966 13662 16966 0 clk_divider.count_out\[27\]
rlabel metal2 24886 9146 24886 9146 0 clk_divider.count_out\[2\]
rlabel metal2 24794 8262 24794 8262 0 clk_divider.count_out\[3\]
rlabel metal2 13938 7327 13938 7327 0 clk_divider.count_out\[4\]
rlabel metal1 13708 7310 13708 7310 0 clk_divider.count_out\[5\]
rlabel metal2 13018 10183 13018 10183 0 clk_divider.count_out\[6\]
rlabel metal2 12834 13498 12834 13498 0 clk_divider.count_out\[7\]
rlabel metal1 13018 12852 13018 12852 0 clk_divider.count_out\[8\]
rlabel metal2 15410 13260 15410 13260 0 clk_divider.count_out\[9\]
rlabel metal1 24380 11322 24380 11322 0 clk_divider.next_count\[0\]
rlabel metal1 16790 11186 16790 11186 0 clk_divider.next_count\[10\]
rlabel metal1 17112 7242 17112 7242 0 clk_divider.next_count\[11\]
rlabel metal1 18262 13770 18262 13770 0 clk_divider.next_count\[12\]
rlabel metal1 18988 6970 18988 6970 0 clk_divider.next_count\[13\]
rlabel metal1 20562 10098 20562 10098 0 clk_divider.next_count\[14\]
rlabel metal1 19780 13226 19780 13226 0 clk_divider.next_count\[15\]
rlabel metal1 23368 13770 23368 13770 0 clk_divider.next_count\[16\]
rlabel metal1 24058 16626 24058 16626 0 clk_divider.next_count\[17\]
rlabel metal1 24150 17782 24150 17782 0 clk_divider.next_count\[18\]
rlabel metal2 17986 17374 17986 17374 0 clk_divider.next_count\[19\]
rlabel metal1 25254 10098 25254 10098 0 clk_divider.next_count\[1\]
rlabel metal1 22540 20026 22540 20026 0 clk_divider.next_count\[20\]
rlabel metal2 19550 20638 19550 20638 0 clk_divider.next_count\[21\]
rlabel metal2 18998 23970 18998 23970 0 clk_divider.next_count\[22\]
rlabel metal1 15824 20570 15824 20570 0 clk_divider.next_count\[23\]
rlabel metal1 11408 20570 11408 20570 0 clk_divider.next_count\[24\]
rlabel metal1 12558 17612 12558 17612 0 clk_divider.next_count\[25\]
rlabel metal1 14950 17544 14950 17544 0 clk_divider.next_count\[26\]
rlabel metal2 13478 17204 13478 17204 0 clk_divider.next_count\[27\]
rlabel metal2 23966 8670 23966 8670 0 clk_divider.next_count\[2\]
rlabel metal2 23782 7582 23782 7582 0 clk_divider.next_count\[3\]
rlabel metal1 15962 7990 15962 7990 0 clk_divider.next_count\[4\]
rlabel metal2 11914 6630 11914 6630 0 clk_divider.next_count\[5\]
rlabel metal2 12466 8126 12466 8126 0 clk_divider.next_count\[6\]
rlabel metal1 11868 13974 11868 13974 0 clk_divider.next_count\[7\]
rlabel metal1 12604 13362 12604 13362 0 clk_divider.next_count\[8\]
rlabel metal2 14674 14110 14674 14110 0 clk_divider.next_count\[9\]
rlabel metal2 21942 17748 21942 17748 0 clk_divider.next_flag
rlabel metal1 24886 21488 24886 21488 0 clk_divider.rollover_flag
rlabel metal1 19320 15878 19320 15878 0 clknet_0_clk
rlabel metal1 14398 13974 14398 13974 0 clknet_2_0__leaf_clk
rlabel metal1 23736 13906 23736 13906 0 clknet_2_1__leaf_clk
rlabel metal1 10672 19890 10672 19890 0 clknet_2_2__leaf_clk
rlabel metal2 26174 17170 26174 17170 0 clknet_2_3__leaf_clk
rlabel metal1 26128 21930 26128 21930 0 count\[0\]
rlabel metal1 27278 20026 27278 20026 0 count\[1\]
rlabel metal1 24472 24718 24472 24718 0 count\[2\]
rlabel metal1 24656 23562 24656 23562 0 count\[3\]
rlabel metal2 23690 23630 23690 23630 0 count\[4\]
rlabel metal1 26082 22950 26082 22950 0 count\[5\]
rlabel metal2 25070 21488 25070 21488 0 counter_to_35.next_count\[0\]
rlabel metal1 25346 20570 25346 20570 0 counter_to_35.next_count\[1\]
rlabel metal1 22218 24582 22218 24582 0 counter_to_35.next_count\[2\]
rlabel via1 22034 23749 22034 23749 0 counter_to_35.next_count\[3\]
rlabel metal1 22356 23290 22356 23290 0 counter_to_35.next_count\[4\]
rlabel metal1 24426 23018 24426 23018 0 counter_to_35.next_count\[5\]
rlabel metal2 25254 19720 25254 19720 0 counter_to_35.next_flag
rlabel metal2 27646 19295 27646 19295 0 done
rlabel metal2 27830 6239 27830 6239 0 enable
rlabel metal2 27646 7106 27646 7106 0 net1
rlabel metal2 2714 13566 2714 13566 0 net10
rlabel metal1 9706 11764 9706 11764 0 net11
rlabel metal2 2622 19652 2622 19652 0 net12
rlabel metal2 2714 20672 2714 20672 0 net13
rlabel metal2 2530 21148 2530 21148 0 net14
rlabel metal1 2208 12818 2208 12818 0 net15
rlabel metal2 1610 19720 1610 19720 0 net16
rlabel metal1 25760 21522 25760 21522 0 net17
rlabel metal2 27830 19142 27830 19142 0 net18
rlabel metal1 23276 27098 23276 27098 0 net19
rlabel metal1 26404 7854 26404 7854 0 net2
rlabel metal1 23874 27642 23874 27642 0 net20
rlabel metal2 25438 27506 25438 27506 0 net21
rlabel metal2 18630 27812 18630 27812 0 net22
rlabel metal1 19182 27302 19182 27302 0 net23
rlabel metal1 16468 28118 16468 28118 0 net24
rlabel metal2 21482 28016 21482 28016 0 net25
rlabel metal1 22356 27642 22356 27642 0 net26
rlabel metal1 22540 27098 22540 27098 0 net27
rlabel metal2 17434 27778 17434 27778 0 net28
rlabel metal2 26818 28084 26818 28084 0 net29
rlabel metal2 15594 7140 15594 7140 0 net3
rlabel metal1 27416 24786 27416 24786 0 net30
rlabel metal2 16974 28050 16974 28050 0 net31
rlabel metal2 21390 28084 21390 28084 0 net32
rlabel metal2 19918 28084 19918 28084 0 net33
rlabel metal1 25438 27098 25438 27098 0 net34
rlabel metal2 17894 27676 17894 27676 0 net35
rlabel metal1 26036 27098 26036 27098 0 net36
rlabel metal1 27094 26010 27094 26010 0 net37
rlabel metal2 24978 28356 24978 28356 0 net38
rlabel metal2 18170 27880 18170 27880 0 net39
rlabel metal1 9982 27472 9982 27472 0 net4
rlabel metal1 18078 28186 18078 28186 0 net40
rlabel metal1 19090 27098 19090 27098 0 net41
rlabel metal1 27554 25296 27554 25296 0 net42
rlabel metal1 27508 24174 27508 24174 0 net43
rlabel metal1 27186 23290 27186 23290 0 net44
rlabel metal1 27462 22610 27462 22610 0 net45
rlabel metal1 27232 27642 27232 27642 0 net46
rlabel metal2 17250 27982 17250 27982 0 net47
rlabel metal1 19642 28186 19642 28186 0 net48
rlabel metal2 17986 27948 17986 27948 0 net49
rlabel metal1 2990 22440 2990 22440 0 net5
rlabel metal1 24426 27642 24426 27642 0 net50
rlabel metal2 20470 28356 20470 28356 0 net51
rlabel metal2 26174 27642 26174 27642 0 net52
rlabel metal1 22770 19754 22770 19754 0 net53
rlabel metal2 22310 14195 22310 14195 0 net54
rlabel metal1 17572 12682 17572 12682 0 net55
rlabel metal2 24012 19244 24012 19244 0 net56
rlabel metal1 12880 18394 12880 18394 0 net57
rlabel metal2 21068 7378 21068 7378 0 net58
rlabel metal1 13938 13158 13938 13158 0 net59
rlabel metal2 1610 23936 1610 23936 0 net6
rlabel via2 24610 13277 24610 13277 0 net60
rlabel metal1 22678 19822 22678 19822 0 net61
rlabel metal1 20976 7378 20976 7378 0 net62
rlabel metal1 20378 14246 20378 14246 0 net63
rlabel metal2 22770 21148 22770 21148 0 net64
rlabel metal1 23920 17646 23920 17646 0 net65
rlabel metal2 21482 26724 21482 26724 0 net66
rlabel metal1 22172 25262 22172 25262 0 net67
rlabel metal1 22034 28016 22034 28016 0 net68
rlabel via1 24242 26554 24242 26554 0 net69
rlabel metal1 2208 21862 2208 21862 0 net7
rlabel metal1 22816 28050 22816 28050 0 net70
rlabel via1 25337 27506 25337 27506 0 net71
rlabel metal2 27002 20944 27002 20944 0 net72
rlabel metal1 25990 21896 25990 21896 0 net73
rlabel metal1 24886 21590 24886 21590 0 net74
rlabel metal2 18446 7684 18446 7684 0 net75
rlabel metal2 21390 20740 21390 20740 0 net76
rlabel metal1 23276 17714 23276 17714 0 net77
rlabel metal1 6486 12206 6486 12206 0 net78
rlabel metal1 6716 27438 6716 27438 0 net79
rlabel metal1 12650 7888 12650 7888 0 net8
rlabel metal1 2438 23732 2438 23732 0 net80
rlabel metal1 12650 25296 12650 25296 0 net81
rlabel metal1 13478 26418 13478 26418 0 net82
rlabel metal1 16245 13974 16245 13974 0 net83
rlabel metal2 25162 13974 25162 13974 0 net84
rlabel metal1 23690 20325 23690 20325 0 net85
rlabel metal3 25231 17204 25231 17204 0 net86
rlabel metal1 2300 17850 2300 17850 0 net87
rlabel metal1 13432 13906 13432 13906 0 net88
rlabel metal2 22310 7599 22310 7599 0 net89
rlabel metal2 1978 10812 1978 10812 0 net9
rlabel metal1 18998 16558 18998 16558 0 net90
rlabel metal1 22310 19720 22310 19720 0 net91
rlabel metal2 27830 5593 27830 5593 0 nrst
rlabel metal1 23460 28730 23460 28730 0 out[0]
rlabel metal2 24150 29767 24150 29767 0 out[10]
rlabel metal1 28244 28186 28244 28186 0 out[11]
rlabel metal2 11822 29767 11822 29767 0 out[12]
rlabel metal2 15686 29767 15686 29767 0 out[13]
rlabel metal2 13110 29767 13110 29767 0 out[14]
rlabel metal2 18262 29767 18262 29767 0 out[15]
rlabel metal2 22034 29767 22034 29767 0 out[16]
rlabel metal2 22862 29767 22862 29767 0 out[17]
rlabel metal2 15042 29767 15042 29767 0 out[18]
rlabel metal2 27370 29767 27370 29767 0 out[19]
rlabel via2 27738 24565 27738 24565 0 out[1]
rlabel metal2 16330 29767 16330 29767 0 out[20]
rlabel metal2 21574 29767 21574 29767 0 out[21]
rlabel metal2 20286 29767 20286 29767 0 out[22]
rlabel metal2 26082 29767 26082 29767 0 out[23]
rlabel metal2 17618 29767 17618 29767 0 out[24]
rlabel metal2 26726 29767 26726 29767 0 out[25]
rlabel metal2 27738 26197 27738 26197 0 out[26]
rlabel metal2 25438 29767 25438 29767 0 out[27]
rlabel metal2 14398 29767 14398 29767 0 out[28]
rlabel metal2 16974 29767 16974 29767 0 out[29]
rlabel metal2 19642 29767 19642 29767 0 out[2]
rlabel metal2 27738 25177 27738 25177 0 out[30]
rlabel metal2 27738 23953 27738 23953 0 out[31]
rlabel metal2 27738 23341 27738 23341 0 out[32]
rlabel via2 27738 22491 27738 22491 0 out[33]
rlabel metal1 27692 27914 27692 27914 0 out[3]
rlabel metal2 12374 29767 12374 29767 0 out[4]
rlabel metal2 18906 29767 18906 29767 0 out[5]
rlabel metal2 13754 29767 13754 29767 0 out[6]
rlabel metal2 24794 29767 24794 29767 0 out[7]
rlabel metal1 20746 28730 20746 28730 0 out[8]
rlabel metal1 27784 28730 27784 28730 0 out[9]
rlabel metal2 9062 1588 9062 1588 0 prescaler[0]
rlabel metal3 1096 23188 1096 23188 0 prescaler[10]
rlabel metal3 751 22508 751 22508 0 prescaler[11]
rlabel metal3 751 23868 751 23868 0 prescaler[12]
rlabel metal3 751 21828 751 21828 0 prescaler[13]
rlabel metal2 5842 1588 5842 1588 0 prescaler[1]
rlabel metal3 751 11628 751 11628 0 prescaler[2]
rlabel metal3 1050 13668 1050 13668 0 prescaler[3]
rlabel metal3 1050 15028 1050 15028 0 prescaler[4]
rlabel metal3 751 17068 751 17068 0 prescaler[5]
rlabel metal3 751 19788 751 19788 0 prescaler[6]
rlabel metal3 866 21148 866 21148 0 prescaler[7]
rlabel metal3 1096 20468 1096 20468 0 prescaler[8]
rlabel metal3 1050 19108 1050 19108 0 prescaler[9]
rlabel via2 27830 14365 27830 14365 0 stop
<< properties >>
string FIXED_BBOX 0 0 29332 31476
<< end >>
